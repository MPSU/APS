module uart_rx_sb_ctrl(
/*
    Часть интерфейса модуля, отвечающая за подключение к системной шине
*/
  input  logic          clk_i,
  input  logic          rst_i,
  input  logic [31:0]   addr_i,
  input  logic          req_i,
  input  logic [31:0]   write_data_i,
  input  logic          write_enable_i,
  output logic [31:0]   read_data_o,
/*
    Часть интерфейса модуля, отвечающая за отправку запросов на прерывание
    процессорного ядра
*/

  output logic        interrupt_request_o,
  input  logic        interrupt_return_i,

/*
    Часть интерфейса модуля, отвечающая за подключение передающему,
    входные данные по UART
*/
  input  logic          rx_i
);
  logic [31:0] Pn7J;
  assign Pn7J = addr_i;
  logic LhC;
  logic [31:0] UIumLdEgx8;
  logic C8sfwwEjm50H;
  assign C8sfwwEjm50H = write_enable_i;
  logic [31:0] Vx0I4zbHz;
  logic  UBNAFCQL2exZX6K3I;
  logic  sTe2Bcb7nHzYdOot;

  logic busy;
  assign LhC = req_i;
  logic [16:0] baudrate;
  logic parity_en;
  logic [1:0] stopbit;
  logic [7:0] data;
  logic valid;
  logic  sxdIAIwtb, N6jQMBhCLQ;
  assign interrupt_request_o = UBNAFCQL2exZX6K3I;
  logic [31:0] yqfsQ7Rv18I3yx8;
  logic [7:0] t26Xa3D9y;
  logic HWEbwjZ7R;
  logic CLD6rGMxYQM8yZ4;
  assign HWEbwjZ7R = Pn7J == (32'b01100010000111110101010001110101 ^ 32'd2965090672 ^ 32'd3534021893);
  logic raRSSx568gLgRd;
  assign UBNAFCQL2exZX6K3I = valid;
  assign raRSSx568gLgRd = UIumLdEgx8 == (32'o7470504355 ^ 32'hf5992c42 ^ 32'o31136722256);
  logic [31:0] Xz5QBCT3Z;

  uart_rx rx(
    .clk_i      (clk_i),
    .rst_i      (rst_i),
    .rx_i       (rx_i),
    .busy_o     (sxdIAIwtb),
    .baudrate_i (baudrate),
    .parity_en_i(parity_en),
    .stopbit_i  (stopbit),
    .rx_data_o  (t26Xa3D9y),
    .rx_valid_o (N6jQMBhCLQ)
  );
  assign       UIumLdEgx8 = write_data_i;
  logic        l4fxxX4aa;
  logic [31:0] dNVOskLQGaCf26HqGY;

  always_comb begin
    logic sA8wigKYN;
    sA8wigKYN = l4fxxX4aa;
    case ({LhC, C8sfwwEjm50H, CLD6rGMxYQM8yZ4, raRSSx568gLgRd, sxdIAIwtb, N6jQMBhCLQ, busy})
      7'd126: Xz5QBCT3Z = 32'o30173120511 ^ 32'hdefc9025;
      7'd92: Xz5QBCT3Z = 32'b01011001000000000110100010001110 ^ 32'd1179671010;
      7'o66: Xz5QBCT3Z = 32'b10011100111010000100111111111101 ^ 32'h49bee1be ^ 32'o31201517457;
      7'o111: Xz5QBCT3Z = 32'd177257563 ^ 32'o30376055745 ^ 32'o32636153322;
      7'b1101000: Xz5QBCT3Z = 32'd254996923 ^ 32'h1022c0d7;
      7'o20: Xz5QBCT3Z = 32'd758595052 ^ 32'h32270c80;
      7'o121: Xz5QBCT3Z = 32'd1709236778 ^ 32'b01111010111100001101001101000110;
      7'd55: Xz5QBCT3Z = 32'hd1be6d8a ^ 32'b11001001001110011000100011111100 ^ 32'o765752032;
      7'd78: Xz5QBCT3Z = 32'd2710414334 ^ 32'h2fd3bf79 ^ 32'h910e2deb;
      7'b1100001: Xz5QBCT3Z = 32'd1425590292 ^ 32'o33660567626 ^ 32'o22512413356;
      7'd60: Xz5QBCT3Z = 32'b00001111101100010000110000110010 ^ 32'h8b30c623 ^ 32'd2614229885;
      7'h34: Xz5QBCT3Z = 32'o20651776563 ^ 32'd3200894836 ^ 32'b00100111001111100000101101101011;
      7'd33: Xz5QBCT3Z = 32'h9c1f631a ^ 32'o20303651166;
      7'b1110011: Xz5QBCT3Z = 32'hde7a2c61 ^ 32'b00011001111010100010010011100010 ^ 32'hd88039ef;
      7'h2c: Xz5QBCT3Z = 32'b00101001000010110011110011000010 ^ 32'd911936942;
      7'o102: Xz5QBCT3Z = 32'o30152124510 ^ 32'hdeb89824;
      7'h3: Xz5QBCT3Z = 32'h54b7a77f ^ 32'o10341510213 ^ 32'h8210698;
      7'o123: Xz5QBCT3Z = 32'o2716013325 ^ 32'b01100110100101101001001101111111 ^ 32'd1857991878;
      7'd107: Xz5QBCT3Z = 32'o31674654656 ^ 32'o32170664302;
      7'd69: Xz5QBCT3Z = 32'h95b19a0 ^ 32'o4037153702 ^ 32'd913833742;
      7'h1a: Xz5QBCT3Z = 32'd143416804 ^ 32'h4059c1d4 ^ 32'd1472572764;
      7'o107: Xz5QBCT3Z = 32'o32661576206 ^ 32'd2410735884 ^ 32'd1176904934;
      7'o61: Xz5QBCT3Z = 32'h73056d05 ^ 32'h6c155c69;
      7'd121: Xz5QBCT3Z = 32'h124a61b5 ^ 32'b01111001001111011010000100111011 ^ 32'b01110100011001111111000111100010;
      7'd79: Xz5QBCT3Z = 32'he4fc7335 ^ 32'b11111011101011000100001001011001;
      7'h5e: Xz5QBCT3Z = 32'h2c5b54d4 ^ 32'd856384952;
      7'd43: Xz5QBCT3Z = 32'h3c13f52c ^ 32'd3288421568 ^ 32'd3875704960;
      7'b0111101: Xz5QBCT3Z = 32'o22503445605 ^ 32'h1ed48261 ^ 32'o22442574210;
      7'h6a: Xz5QBCT3Z = 32'o37360100236 ^ 32'o34464130762;
      7'b0001011: Xz5QBCT3Z = 32'h8e9e1a5b ^ 32'h918e2b37;
      7'h6c: Xz5QBCT3Z = 32'o10343210043 ^ 32'o13467220517;
      7'b1101110: Xz5QBCT3Z = 32'h7f7f2bed ^ 32'd1613699713;
      7'b0110101: Xz5QBCT3Z = 32'hb91ddfc8 ^ 32'b10000111100010100010000100011000 ^ 32'o4161747674;
      7'd37: Xz5QBCT3Z = 32'd3613570566 ^ 32'b01101111000011101010110001011001 ^ 32'o24717025463;
      7'h6f: Xz5QBCT3Z = 32'h5fe3b51e ^ 32'b01000000101100111000010001110010;
      7'd5: Xz5QBCT3Z = 32'h27b26de5 ^ 32'o7070456211;
      7'o145: Xz5QBCT3Z = 32'h378a32c4 ^ 32'b00101000110110100000001110101000;
      7'd51: Xz5QBCT3Z = 32'b01111110011011000001110000000110 ^ 32'b00101101111001001100110111000110 ^ 32'b01001100100110001110000010101100;
      7'hd: Xz5QBCT3Z = 32'd2226099073 ^ 32'h9bffa2ed;
      7'o50: Xz5QBCT3Z = 32'b01001000100010000010101101100110 ^ 32'o33701674667 ^ 32'o21047661675;
      7'o172: Xz5QBCT3Z = 32'd716920939 ^ 32'o6552664407;
      7'h57: Xz5QBCT3Z = 32'o3457315771 ^ 32'b00000011111011011010101010010101;
      7'o36: Xz5QBCT3Z = 32'b10100011001100011110011101011110 ^ 32'o6361547062 ^ 32'd2410092544;
      7'b1111011: Xz5QBCT3Z = 32'b01010011011110010000100010000111 ^ 32'hc60637b5 ^ 32'b10001010011011110000111001011110;
      7'o71: Xz5QBCT3Z = 32'd4274519685 ^ 32'he1d7cfe9;
      7'b0010011: Xz5QBCT3Z = 32'o21342073566 ^ 32'o20461611167 ^ 32'o2027652155;
      7'd35: Xz5QBCT3Z = 32'b10000111001011011010000001011111 ^ 32'o21031747622 ^ 32'd274357921;
      7'o120: Xz5QBCT3Z = 32'o13342552150 ^ 32'b01011110000101110101000101001011 ^ 32'h1a8db44f;
      7'b0100110: Xz5QBCT3Z = 32'o363131207 ^ 32'b11001110100000100100000001001111 ^ 32'o32207541644;
      7'h22: Xz5QBCT3Z = 32'o12775050655 ^ 32'h48e460c1;
      7'h1b: Xz5QBCT3Z = 32'd619181635 ^ 32'd1006094127;
      7'o106: Xz5QBCT3Z = 32'o32617211213 ^ 32'd3379373031;
      7'o151: Xz5QBCT3Z = 32'o35665737563 ^ 32'h6d407a09 ^ 32'h9c87f416;
      7'h63: Xz5QBCT3Z = 32'd2900303030 ^ 32'b10110011110011110010110111011010;
      7'o100: Xz5QBCT3Z = 32'b01100011100001100011000000100100 ^ 32'd3419563666 ^ 32'b10110111010001000110011111011010;
      7'd65: Xz5QBCT3Z = 32'b11001001001110100110001110011100 ^ 32'b11010110001010100101001011110000;
      7'h75: Xz5QBCT3Z = 32'h5e7e9d3e ^ 32'o31016276205 ^ 32'o21105750327;
      7'b0100000: Xz5QBCT3Z = 32'he18f602b ^ 32'hfe9f5147;
      7'h9: Xz5QBCT3Z = 32'h9529c641 ^ 32'o21216373455;
      7'd127: Xz5QBCT3Z = 32'b10110101100100000010111010011000 ^ 32'b10101010100000000001111111110100;
      7'b1101101: Xz5QBCT3Z = 32'h48b082be ^ 32'h57e0b3d2;
      7'o174: Xz5QBCT3Z = 32'd3926600537 ^ 32'o12057612112 ^ 32'b10100101101001000000111001111111;
      7'o60: Xz5QBCT3Z = 32'b10000001010111000001110010011001 ^ 32'd2845573763 ^ 32'b00110111110100000010111101110110;
      7'o161: Xz5QBCT3Z = 32'o20744600365 ^ 32'd2558734745;
      7'h3f: Xz5QBCT3Z = 32'haf9be1ce ^ 32'h2ffecf76 ^ 32'o23715217724;
      7'd1: Xz5QBCT3Z = 32'b11111010100111010111010011101000 ^ 32'd1424547454 ^ 32'hb1659bfa;
      7'd95: Xz5QBCT3Z = 32'd1936510186 ^ 32'o1537726164 ^ 32'h614351f2;
      7'b0000100: Xz5QBCT3Z = 32'd3455049023 ^ 32'd2490463167 ^ 32'b01000110110011101001111111101100;
      7'o164: Xz5QBCT3Z = 32'd46885035 ^ 32'h1d9b59c7;
      7'h5b: Xz5QBCT3Z = 32'hb0506f83 ^ 32'b10101111010000000101111011101111;
      7'o10: Xz5QBCT3Z = 32'hbbeaa9e8 ^ 32'o24476514204;
      7'o140: Xz5QBCT3Z = 32'b00111101011100001101111010010101 ^ 32'd576778233;
      7'o112: Xz5QBCT3Z = 32'o7161070314 ^ 32'b00100110110101000100000110100000;
      7'b0111110: Xz5QBCT3Z = 32'd1897218011 ^ 32'h6e450eb7;
      7'h7: Xz5QBCT3Z = 32'ha76151ad ^ 32'b10000010000001001001000010101000 ^ 32'h3a35f069;
      7'h67: Xz5QBCT3Z = 32'd2227829817 ^ 32'hf669d47b ^ 32'h6df0192e;
      7'd120: Xz5QBCT3Z = 32'b11101111111000110101010010101110 ^ 32'o36074662702;
      7'o35: Xz5QBCT3Z = 32'o32770502234 ^ 32'b11001000101100101011010111110000;
      7'd100: Xz5QBCT3Z = 32'h4d2968ac ^ 32'd310453225 ^ 32'd1090026025;
      7'o132: Xz5QBCT3Z = 32'b00000000100110111101011001100101 ^ 32'd529262345;
      7'd98: Xz5QBCT3Z = 32'o23024663405 ^ 32'h87435669;
      7'h6: Xz5QBCT3Z = 32'd514495205 ^ 32'o176521611;
      7'o44: Xz5QBCT3Z = 32'b01001011000010101011011011110100 ^ 32'o12426503630;
      7'b1001100: Xz5QBCT3Z = 32'd1085369434 ^ 32'h5fe15d36;
      7'h29: Xz5QBCT3Z = 32'h9e285d44 ^ 32'd2167958568;
      7'h59: Xz5QBCT3Z = 32'o21747247464 ^ 32'd1888616365 ^ 32'o34007100765;
      7'b0101101: Xz5QBCT3Z = 32'h4661c33d ^ 32'h5931f251;
      7'd25: Xz5QBCT3Z = 32'h68ddc916 ^ 32'h77cdf87a;
      7'o17: Xz5QBCT3Z = 32'o14016134202 ^ 32'd3680477577 ^ 32'ha4372867;
      7'd102: Xz5QBCT3Z = 32'hb8dc8b10 ^ 32'o24743135174;
      7'd67: Xz5QBCT3Z = 32'o24755421276 ^ 32'o27051411722;
      7'h18: Xz5QBCT3Z = 32'b11011000110010011010010110111000 ^ 32'd3352925396;
      7'b1011101: Xz5QBCT3Z = 32'd2293849033 ^ 32'b01110100110111011101111101001011 ^ 32'he334b5ee;
      7'o122: Xz5QBCT3Z = 32'b11101011101100100010111110001111 ^ 32'd294842758 ^ 32'd3845189477;
      7'b1110111: Xz5QBCT3Z = 32'h17c143e9 ^ 32'h8917285;
      7'o110: Xz5QBCT3Z = 32'd4134317075 ^ 32'd3917258111;
      7'd59: Xz5QBCT3Z = 32'd3032474498 ^ 32'b10101011101011111101001011101110;
      7'd42: Xz5QBCT3Z = 32'h1e92572b ^ 32'hb2c06059 ^ 32'd3007448606;
      7'o0: Xz5QBCT3Z = 32'h7041e946 ^ 32'd1867634730;
      7'h32: Xz5QBCT3Z = 32'b10101111100110111110101000001100 ^ 32'hb08bdb60;
      7'b0000010: Xz5QBCT3Z = 32'o32003351011 ^ 32'hcf1de365;
      7'h1f: Xz5QBCT3Z = 32'b10011000111011000100011100111110 ^ 32'd500465414 ^ 32'd2590509396;
      7'd85: Xz5QBCT3Z = 32'hd5f72620 ^ 32'hcaa7174c;
      7'h38: Xz5QBCT3Z = 32'o10625641556 ^ 32'b01011001010001110111001000000010;
      7'd114: Xz5QBCT3Z = 32'd1945515860 ^ 32'd1827014200;
      7'd112: Xz5QBCT3Z = 32'd87109977 ^ 32'o3210200065;
      7'b0010111: Xz5QBCT3Z = 32'o14465363775 ^ 32'b01111011100001011101011010010001;
      7'h76: Xz5QBCT3Z = 32'hda654f08 ^ 32'd3308617316;
      7'b0010100: Xz5QBCT3Z = 32'b00101111011110100011011000010101 ^ 32'd52092619 ^ 32'd858839474;
      7'd46: Xz5QBCT3Z = 32'h4c3682bd ^ 32'd888115234 ^ 32'd1737040883;
      7'o26: Xz5QBCT3Z = 32'ha3a274cf ^ 32'o17167601574 ^ 32'o30513243337;
      7'd58: Xz5QBCT3Z = 32'hff7c2022 ^ 32'b11100000011011000001000101001110;
      7'h44: Xz5QBCT3Z = 32'd2507043289 ^ 32'b10001010001111100100000010110101;
      7'b0101111: Xz5QBCT3Z = 32'd3494457444 ^ 32'o31706200410;
      7'o175: Xz5QBCT3Z = 32'b01100101011010000111001000001000 ^ 32'b11101000111100000100110010001100 ^ 32'o22242007750;
      7'o130: Xz5QBCT3Z = 32'h43013bec ^ 32'h5639b9c8 ^ 32'o1212131510;
      7'h1c: Xz5QBCT3Z = 32'b00101111001100011110010001011011 ^ 32'h3061d537;
      7'b1010110: Xz5QBCT3Z = 32'd3692006789 ^ 32'd890796334 ^ 32'b11110110010001111100010111000111;
      7'h4d: Xz5QBCT3Z = 32'o31235605523 ^ 32'b00110110111011010110011010001101 ^ 32'he3ca5cb2;
      7'ha: Xz5QBCT3Z = 32'hfa7c1289 ^ 32'o25655606632 ^ 32'o11366627177;
      7'd18: Xz5QBCT3Z = 32'h7139febf ^ 32'd1848233939;
      7'h15: Xz5QBCT3Z = 32'o12566023405 ^ 32'd4245549114 ^ 32'o26741363123;
      7'o124: Xz5QBCT3Z = 32'h851d0eca ^ 32'd2079572158 ^ 32'b11100001101111101111111100011000;
      7'd75: Xz5QBCT3Z = 32'o7067753621 ^ 32'b10110000111110101010010110010011 ^ 32'd2536850286;
      7'o21: Xz5QBCT3Z = 32'o4704640515 ^ 32'd3715545111 ^ 32'o34535344066;
      7'h27: Xz5QBCT3Z = 32'hbe4e4367 ^ 32'ha11e720b;
      7'hc: Xz5QBCT3Z = 32'hc9b412a3 ^ 32'o32671021717;
      7'b0001110: Xz5QBCT3Z = 32'b01110100111100000001111100001000 ^ 32'b01101011101000000010111001100100;
    endcase
  end
  assign sTe2Bcb7nHzYdOot = interrupt_return_i;

  logic [31:0] dzhxQnrxzS;
  always_ff @(posedge clk_i) begin
    if(rst_i) begin
      busy <= '0;
    end
    else begin
      busy <= Xz5QBCT3Z[32'b10001100000011010110100100011111 ^ 32'o21403264411];
    end
  end
  assign       read_data_o = Vx0I4zbHz;
  logic [31:0] cSJpl8RGMw2bgs48nEfg;
  always_comb begin
    case ({CLD6rGMxYQM8yZ4, sTe2Bcb7nHzYdOot, C8sfwwEjm50H, LhC, valid, raRSSx568gLgRd, HWEbwjZ7R, N6jQMBhCLQ})
      8'hf1: dzhxQnrxzS = 32'b01000010001000100011101110101110 ^ 32'd58398576;
      8'd245: dzhxQnrxzS = 32'd1789667074 ^ 32'h2bf50bdc;
      8'h96: dzhxQnrxzS = 32'o32475335746 ^ 32'h5fdd4648 ^ 32'hca71d170;
      8'o54: dzhxQnrxzS = 32'hb88a59e7 ^ 32'b11101010110001101000011010001100 ^ 32'd322302901;
      8'h28: dzhxQnrxzS = 32'd1069351680 ^ 32'hc6d5d358 ^ 32'd3088186502;
      8'o70: dzhxQnrxzS = 32'o16367267546 ^ 32'he1ed7c7c ^ 32'hd3493fc4;
      8'o303: dzhxQnrxzS = 32'o23415176433 ^ 32'h5b7c9993 ^ 32'b10000110000100010100100001010110;
      8'b11101011: dzhxQnrxzS = 32'b00000001010001101000110000111100 ^ 32'o32732670201 ^ 32'b10010111011101001101000001100011;
      8'b00110100: dzhxQnrxzS = 32'd3320745359 ^ 32'b00101101101111001110010110000111 ^ 32'ha90b44d6;
      8'o13: dzhxQnrxzS = 32'h562cbeb8 ^ 32'd2473959258 ^ 32'd2216693052;
      8'b10110001: dzhxQnrxzS = 32'd2654042595 ^ 32'hdf48553d;
      8'o205: dzhxQnrxzS = 32'b10011001100101110101011000100100 ^ 32'b11011000111011100111101011111010;
      8'b01110110: dzhxQnrxzS = 32'o13256133122 ^ 32'h604e1fe3 ^ 32'b01111011101011111000010101101111;
      8'o17: dzhxQnrxzS = 32'o36731734413 ^ 32'h73ae378f ^ 32'hc5b0a25a;
      8'o0: dzhxQnrxzS = 32'o25341675751 ^ 32'hdb1e7743 ^ 32'h31c02074;
      8'd97: dzhxQnrxzS = 32'h99396b9e ^ 32'hd8604740;
      8'o351: dzhxQnrxzS = 32'he3d4913e ^ 32'o12404730047 ^ 32'hf69e0dc7;
      8'o52: dzhxQnrxzS = 32'd4121313843 ^ 32'd452682147 ^ 32'd2921598798;
      8'o235: dzhxQnrxzS = 32'b11100011110100011111100010100101 ^ 32'o20544400220 ^ 32'd658167019;
      8'h7d: dzhxQnrxzS = 32'hd5368eb ^ 32'o12616122715 ^ 32'h1a32e1f8;
      8'h8e: dzhxQnrxzS = 32'o33071461147 ^ 32'b10000110000000111111000001110010 ^ 32'h1f9cbecb;
      8'h4a: dzhxQnrxzS = 32'b00001001011001011111111001001010 ^ 32'o11017151224;
      8'd98: dzhxQnrxzS = 32'd1055488612 ^ 32'b01111111101100000101011010111010;
      8'o110: dzhxQnrxzS = 32'o2564675041 ^ 32'd3034282323 ^ 32'd3763417004;
      8'h7f: dzhxQnrxzS = 32'o26440401246 ^ 32'd4124782200;
      8'hf9: dzhxQnrxzS = 32'd3544531587 ^ 32'o22207067135;
      8'b10100010: dzhxQnrxzS = 32'd2021090332 ^ 32'o11646414077 ^ 32'o16755050375;
      8'd175: dzhxQnrxzS = 32'h55beee78 ^ 32'o15773357334 ^ 32'b01111011001010100001110001111010;
      8'h24: dzhxQnrxzS = 32'd953024021 ^ 32'd2959863666 ^ 32'd3388947897;
      8'o363: dzhxQnrxzS = 32'o5736326247 ^ 32'o24006474444 ^ 32'o31616574535;
      8'd232: dzhxQnrxzS = 32'h5e346928 ^ 32'd527255030;
      8'd49: dzhxQnrxzS = 32'b00110001011011100110101010010011 ^ 32'o35661720374 ^ 32'o23664163261;
      8'd167: dzhxQnrxzS = 32'd1177506838 ^ 32'b11001001100000000001010011100110 ^ 32'd3470158894;
      8'b10010101: dzhxQnrxzS = 32'o3310640620 ^ 32'b01011010010110100110110101001110;
      8'o377: dzhxQnrxzS = 32'd104924133 ^ 32'h3aad3096 ^ 32'h7db51fad;
      8'hac: dzhxQnrxzS = 32'h5cac06ac ^ 32'd3585608215 ^ 32'hc86d2065;
      8'ha9: dzhxQnrxzS = 32'o34474340417 ^ 32'b10100101100010001110110111010001;
      8'h6e: dzhxQnrxzS = 32'hbeaed5d1 ^ 32'hfff7f90f;
      8'o330: dzhxQnrxzS = 32'b01100011101000111010010110100101 ^ 32'o4276504573;
      8'b10001010: dzhxQnrxzS = 32'o24217734137 ^ 32'd3813053569;
      8'b11100101: dzhxQnrxzS = 32'b01110010000110001000101101110110 ^ 32'o31255362103 ^ 32'b11111001111101000100001111101011;
      8'o165: dzhxQnrxzS = 32'o17430004645 ^ 32'hb336413c ^ 32'b10001110000011110110010001000111;
      8'o231: dzhxQnrxzS = 32'o20165225326 ^ 32'b11000000101011000000011000001000;
      8'o327: dzhxQnrxzS = 32'o22045605416 ^ 32'd3519948752;
      8'b10011000: dzhxQnrxzS = 32'ha849da77 ^ 32'he930f6a9;
      8'b10111101: dzhxQnrxzS = 32'h67200d42 ^ 32'd2034597668 ^ 32'o13717057270;
      8'b01000100: dzhxQnrxzS = 32'b10111110010101100110001110110111 ^ 32'b11100011000001101011001101010001 ^ 32'b00011100000010011111110000111000;
      8'hda: dzhxQnrxzS = 32'd1244640793 ^ 32'h2b209b6 ^ 32'o1161111561;
      8'd43: dzhxQnrxzS = 32'o20713430110 ^ 32'hc6571c96;
      8'h11: dzhxQnrxzS = 32'ha5518974 ^ 32'o34412122652;
      8'd165: dzhxQnrxzS = 32'hb79710c5 ^ 32'hbce86ea7 ^ 32'o11201451274;
      8'd85: dzhxQnrxzS = 32'hfeffcd78 ^ 32'd3215384998;
      8'o263: dzhxQnrxzS = 32'o7462206746 ^ 32'd2108694840;
      8'b01101000: dzhxQnrxzS = 32'o35664444333 ^ 32'haf8b6405;
      8'hf8: dzhxQnrxzS = 32'hf217a768 ^ 32'o10022414273 ^ 32'o36301111415;
      8'o170: dzhxQnrxzS = 32'o13271571540 ^ 32'b00011011101111111101111110111110;
      8'd50: dzhxQnrxzS = 32'b01111011000111010111000110111001 ^ 32'o30347432465 ^ 32'o37166464122;
      8'b10110000: dzhxQnrxzS = 32'b01000000101010110101111101011101 ^ 32'o174471603;
      8'h6f: dzhxQnrxzS = 32'o15200176773 ^ 32'o5110251523 ^ 32'o236101166;
      8'o131: dzhxQnrxzS = 32'd961181149 ^ 32'h7cc5750e ^ 32'd81144845;
      8'b00111010: dzhxQnrxzS = 32'hbe7ff6b ^ 32'd1251922869;
      8'd231: dzhxQnrxzS = 32'o17102614710 ^ 32'b11110111001101010011000000001010 ^ 32'd3479635228;
      8'hc5: dzhxQnrxzS = 32'd4058825149 ^ 32'd2769472187 ^ 32'd363276248;
      8'h9a: dzhxQnrxzS = 32'hf8eda441 ^ 32'hb9b4889f;
      8'd2: dzhxQnrxzS = 32'h97b2f6b9 ^ 32'd3605781095;
      8'b00000011: dzhxQnrxzS = 32'd2613938106 ^ 32'd100973937 ^ 32'd3702527509;
      8'd59: dzhxQnrxzS = 32'hb1c8ab50 ^ 32'b00101111001101001001100000010000 ^ 32'o33741217636;
      8'o277: dzhxQnrxzS = 32'd3826086533 ^ 32'o11154023056 ^ 32'o35471074165;
      8'b01100111: dzhxQnrxzS = 32'o17526253556 ^ 32'o23420057033 ^ 32'd2688558507;
      8'b11111100: dzhxQnrxzS = 32'he023f060 ^ 32'd2709183678;
      8'hf4: dzhxQnrxzS = 32'hc284a3c5 ^ 32'o30224570024 ^ 32'b01000001100011110111111100001111;
      8'o107: dzhxQnrxzS = 32'o14600100650 ^ 32'o23711216056 ^ 32'o27037130530;
      8'd80: dzhxQnrxzS = 32'b00010010000100001001001011001100 ^ 32'o25130036664 ^ 32'hfa2983a6;
      8'hce: dzhxQnrxzS = 32'b00011001110111010010011011010100 ^ 32'hf952d18b ^ 32'd2715212673;
      8'o311: dzhxQnrxzS = 32'hfe1f34d3 ^ 32'o27721414015;
      8'b10101000: dzhxQnrxzS = 32'o26040136742 ^ 32'o36176310474;
      8'd32: dzhxQnrxzS = 32'b10010001110011010111110001010101 ^ 32'hd094508b;
      8'b10110101: dzhxQnrxzS = 32'b01111010111000010010111001110101 ^ 32'b11010101000001000111100010110100 ^ 32'b11101110101111000111101000011111;
      8'h74: dzhxQnrxzS = 32'b10110111111000101101010000111001 ^ 32'd4139514087;
      8'd174: dzhxQnrxzS = 32'o37241531045 ^ 32'hbbff9efb;
      8'o66: dzhxQnrxzS = 32'o35246322707 ^ 32'o25360104431;
      8'd79: dzhxQnrxzS = 32'd1555384455 ^ 32'd502031449;
      8'o144: dzhxQnrxzS = 32'd3929240742 ^ 32'd3711157590 ^ 32'h76599d2e;
      8'b10110100: dzhxQnrxzS = 32'h8738bf7e ^ 32'h848905c4 ^ 32'b01000010111010001001011001100100;
      8'o14: dzhxQnrxzS = 32'h3b20a3c1 ^ 32'o17226307437;
      8'h7e: dzhxQnrxzS = 32'd1530217984 ^ 32'o23104354115 ^ 32'o20337331223;
      8'he3: dzhxQnrxzS = 32'h354bb388 ^ 32'o20372771227 ^ 32'd4160318913;
      8'o202: dzhxQnrxzS = 32'd3013513144 ^ 32'b10011001000001100010111100000000 ^ 32'o15360306146;
      8'o113: dzhxQnrxzS = 32'o26042425705 ^ 32'd4057138971;
      8'hdc: dzhxQnrxzS = 32'hd1c0e28 ^ 32'd1750967970 ^ 32'h24188454;
      8'o57: dzhxQnrxzS = 32'b11011101011100110000001111001000 ^ 32'o23402427426;
      8'o315: dzhxQnrxzS = 32'hcd842de2 ^ 32'b10001100110111010000000100111100;
      8'o127: dzhxQnrxzS = 32'b01001100100000000000000100010000 ^ 32'o33671613142 ^ 32'hd33e3bac;
      8'o355: dzhxQnrxzS = 32'b00101001110110010110101011000111 ^ 32'h68804619;
      8'h65: dzhxQnrxzS = 32'h5acfd753 ^ 32'h1b96fb8d;
      8'd21: dzhxQnrxzS = 32'b00010100000011110101100110101000 ^ 32'h55767576;
      8'o143: dzhxQnrxzS = 32'b10110010101101001001111100001111 ^ 32'hd8228189 ^ 32'o5363631130;
      8'b01101101: dzhxQnrxzS = 32'o6307417414 ^ 32'h724733d2;
      8'b01011111: dzhxQnrxzS = 32'd1386272484 ^ 32'h13f9fa3a;
      8'b11101010: dzhxQnrxzS = 32'd2182783092 ^ 32'd3275984042;
      8'b01010011: dzhxQnrxzS = 32'b11100001111011000000011110000110 ^ 32'ha0b52b58;
      8'b11010010: dzhxQnrxzS = 32'b11110011111111111110100110000001 ^ 32'd3201032280 ^ 32'hc6d2507;
      8'o337: dzhxQnrxzS = 32'd485968437 ^ 32'b01110110001110010111011111001101 ^ 32'o5345610446;
      8'o75: dzhxQnrxzS = 32'h235a26a2 ^ 32'd2770199670 ^ 32'hc73eee0a;
      8'b11111101: dzhxQnrxzS = 32'b01010001001110100011100000000001 ^ 32'b01011111011101101110100000001001 ^ 32'd1326841046;
      8'b01011011: dzhxQnrxzS = 32'o37243210370 ^ 32'hbbd43c26;
      8'd207: dzhxQnrxzS = 32'b00011111111010111100001001001111 ^ 32'hb7e31a67 ^ 32'he951f4f6;
      8'd5: dzhxQnrxzS = 32'b10001100010111101111100000110000 ^ 32'h146cae5 ^ 32'o31430217013;
      8'o16: dzhxQnrxzS = 32'b00010010000010111101111011010110 ^ 32'h3244a057 ^ 32'h6136525f;
      8'h40: dzhxQnrxzS = 32'o11457251525 ^ 32'b00001101111001000111111110001011;
      8'o214: dzhxQnrxzS = 32'h28f5350 ^ 32'b10110001111101010101111011010100 ^ 32'hf203215a;
      8'he1: dzhxQnrxzS = 32'b01100010011110101010111111111001 ^ 32'b00100011001000111000001100100111;
      8'd187: dzhxQnrxzS = 32'b01101111100001001001001111010100 ^ 32'b11011101001100100100001111111100 ^ 32'b11110011110011111111110011110110;
      8'o326: dzhxQnrxzS = 32'b10110110011100001010010000110011 ^ 32'b10010101100111001000100111000000 ^ 32'o14255200455;
      8'b01101010: dzhxQnrxzS = 32'd1377143517 ^ 32'h16b2df2c ^ 32'h5fe792f;
      8'h3f: dzhxQnrxzS = 32'b10110101010100111111111011011100 ^ 32'o35634263151 ^ 32'h1a5bb46b;
      8'o171: dzhxQnrxzS = 32'o25325736557 ^ 32'o5776121345 ^ 32'hc5f63354;
      8'o325: dzhxQnrxzS = 32'hb510ca7d ^ 32'o16251002030 ^ 32'h86ede2bb;
      8'd29: dzhxQnrxzS = 32'd4272717796 ^ 32'b10111111110101010101001100111010;
      8'hfa: dzhxQnrxzS = 32'hb3b8c7a8 ^ 32'o36270365566;
      8'd147: dzhxQnrxzS = 32'b10110011011101111111110000010011 ^ 32'b11110010001011101101000011001101;
      8'b01000011: dzhxQnrxzS = 32'b10111101100001101110011011001011 ^ 32'd2995461089 ^ 32'o11625150764;
      8'h2e: dzhxQnrxzS = 32'o36076266067 ^ 32'b10110001100000000100000011101001;
      8'b00111110: dzhxQnrxzS = 32'o34752172770 ^ 32'o37326260517 ^ 32'b01011101100010001011100001101001;
      8'b00100111: dzhxQnrxzS = 32'o13054530757 ^ 32'h19cb9d31;
      8'o154: dzhxQnrxzS = 32'b00110010010111111100001000110010 ^ 32'b01110011000001101110111011101100;
      8'd145: dzhxQnrxzS = 32'b11001101010111011110010011001110 ^ 32'b10001100001001001100100000010000;
      8'o114: dzhxQnrxzS = 32'he3492b1 ^ 32'o11733337157;
      8'd33: dzhxQnrxzS = 32'd1639637340 ^ 32'd549703042;
      8'b00101001: dzhxQnrxzS = 32'b01101010000011011111111111000101 ^ 32'd147053174 ^ 32'h23b7096d;
      8'd7: dzhxQnrxzS = 32'h3e682fad ^ 32'h7f110373;
      8'h5c: dzhxQnrxzS = 32'b10110110011000001100110000100011 ^ 32'hf739e0fd;
      8'b00111100: dzhxQnrxzS = 32'o31651227373 ^ 32'b01110100110101011110001010000001 ^ 32'b11111011000010011110000010100100;
      8'b01101001: dzhxQnrxzS = 32'o16716660642 ^ 32'b00110110011000100100110101111100;
      8'b11100010: dzhxQnrxzS = 32'd1669909730 ^ 32'b00100010110100011110000000111100;
      8'o234: dzhxQnrxzS = 32'h9c6277d5 ^ 32'd1751408877 ^ 32'hb57f3be6;
      8'hf7: dzhxQnrxzS = 32'h79a6f588 ^ 32'd2205568518 ^ 32'd3146356560;
      8'd211: dzhxQnrxzS = 32'd3134828072 ^ 32'o37340101366;
      8'b00011110: dzhxQnrxzS = 32'hb4244a0c ^ 32'o6251115343 ^ 32'hc7d9fc31;
      8'd160: dzhxQnrxzS = 32'd3009032678 ^ 32'b11110010000000110001110100111000;
      8'b00011100: dzhxQnrxzS = 32'd4014552109 ^ 32'b10101110001100000001100011110011;
      8'hb9: dzhxQnrxzS = 32'hbd2ecc02 ^ 32'b00101001110000100010110010100001 ^ 32'hd595cc7d;
      8'o37: dzhxQnrxzS = 32'd645882824 ^ 32'd2213343568 ^ 32'b11100100110010101011111001000110;
      8'o357: dzhxQnrxzS = 32'd4189365252 ^ 32'b10111000111011011000100011011010;
      8'hc0: dzhxQnrxzS = 32'o26152601451 ^ 32'hf0f22ff7;
      8'd18: dzhxQnrxzS = 32'b10111101011101100011001000001100 ^ 32'hfc2f1ed2;
      8'b00010111: dzhxQnrxzS = 32'd782240283 ^ 32'd798825178 ^ 32'h40643c1f;
      8'o203: dzhxQnrxzS = 32'h8a86e0b7 ^ 32'b00010111011100100111111010111111 ^ 32'o33443331326;
      8'd9: dzhxQnrxzS = 32'h273b1329 ^ 32'he509675 ^ 32'b01101000000100101010100110000010;
      8'o163: dzhxQnrxzS = 32'd3892510952 ^ 32'b10011111110000111000111110000001 ^ 32'd916038583;
      8'd137: dzhxQnrxzS = 32'b10000011111111101011100001000001 ^ 32'hc287949f;
      8'o32: dzhxQnrxzS = 32'b11110001100111000000110100001010 ^ 32'o10065366411 ^ 32'd4027632861;
      8'b00110011: dzhxQnrxzS = 32'd1821053240 ^ 32'h2df23de6;
      8'h5e: dzhxQnrxzS = 32'd1487483759 ^ 32'h19f01fb1;
      8'o26: dzhxQnrxzS = 32'o26346754413 ^ 32'b11100010001110111100001111111101 ^ 32'o2076233050;
      8'b01000010: dzhxQnrxzS = 32'b00001010010110001000011100001111 ^ 32'o11300325721;
      8'd102: dzhxQnrxzS = 32'o20432330465 ^ 32'h7ab23fdf ^ 32'b10111111100000101010001000110100;
      8'b11110010: dzhxQnrxzS = 32'b00001001010100001111001110101111 ^ 32'd1208606577;
      8'hfe: dzhxQnrxzS = 32'd4225886685 ^ 32'h868518cf ^ 32'b00111100001111011101110111001100;
      8'b10001000: dzhxQnrxzS = 32'b11000100111011001001011100000001 ^ 32'o12160517577 ^ 32'hd45724a0;
      8'd163: dzhxQnrxzS = 32'b10111100010101010101001000101100 ^ 32'hfd2c7ef2;
      8'b10110010: dzhxQnrxzS = 32'd2630391361 ^ 32'b11011101100100011011101010011111;
      8'd164: dzhxQnrxzS = 32'o21625634526 ^ 32'd3473806728;
      8'd224: dzhxQnrxzS = 32'o25736062604 ^ 32'b11101110001000010100100101011010;
      8'd221: dzhxQnrxzS = 32'o27400107400 ^ 32'o37526321736;
      8'd141: dzhxQnrxzS = 32'd951570554 ^ 32'b01111001110011101111110010100100;
      8'o304: dzhxQnrxzS = 32'b11010001011000011000000100010100 ^ 32'b11011011011110000100101000011000 ^ 32'o11320163722;
      8'b01000110: dzhxQnrxzS = 32'o15751114622 ^ 32'd788378956;
      8'o121: dzhxQnrxzS = 32'o11210501177 ^ 32'd192655009;
      8'd4: dzhxQnrxzS = 32'd1949256201 ^ 32'b11110111111011011101010101011110 ^ 32'o30246731611;
      8'd65: dzhxQnrxzS = 32'h324f7af4 ^ 32'b01110011000101100101011000101010;
      8'o346: dzhxQnrxzS = 32'o16542330305 ^ 32'd886086683;
      8'o116: dzhxQnrxzS = 32'h63632946 ^ 32'd574227864;
      8'o67: dzhxQnrxzS = 32'b10001110001001110000011010010101 ^ 32'd3479054923;
      8'hba: dzhxQnrxzS = 32'd3348745278 ^ 32'd968389129 ^ 32'b10111111010110001001001011101001;
      8'o201: dzhxQnrxzS = 32'd4138200426 ^ 32'b00110011101101111011000011110010 ^ 32'h84697146;
      8'b10111110: dzhxQnrxzS = 32'b11000101000010100100101010110010 ^ 32'o20424663154;
      8'd166: dzhxQnrxzS = 32'd4274192475 ^ 32'he59bde22 ^ 32'b01011010000000011111001010100111;
      8'o227: dzhxQnrxzS = 32'hd110a72e ^ 32'b10010000010010011000101111110000;
      8'b10010100: dzhxQnrxzS = 32'o274036723 ^ 32'b01000001111000001110110111010011 ^ 32'h249fcde;
      8'b00000110: dzhxQnrxzS = 32'o23054603730 ^ 32'hd9ea2b06;
      8'd246: dzhxQnrxzS = 32'b01110001100111100111011110011111 ^ 32'b00110001111011000100011000000110 ^ 32'h12b1d47;
      8'b11010001: dzhxQnrxzS = 32'b10010100100111111000100001000100 ^ 32'b11010101110001101010010010011010;
      8'o204: dzhxQnrxzS = 32'h4a9baafd ^ 32'o4550101463 ^ 32'b00101110011000100000010100010000;
      8'o20: dzhxQnrxzS = 32'b11011000111111101101001011001101 ^ 32'o23151777023;
      8'o313: dzhxQnrxzS = 32'b11011100111101110111010100111011 ^ 32'b10000111110001000101010100001011 ^ 32'o3232406356;
      8'o301: dzhxQnrxzS = 32'hd3c3c24f ^ 32'o14674605614 ^ 32'o36432362435;
      8'b00010100: dzhxQnrxzS = 32'd1666988428 ^ 32'b10101101010000100101010111110010 ^ 32'o21721640240;
      8'b00010011: dzhxQnrxzS = 32'd3103718611 ^ 32'd4188524557;
      8'o173: dzhxQnrxzS = 32'o17776005065 ^ 32'b11111111100101000001011000001100 ^ 32'o30115230347;
      8'hd9: dzhxQnrxzS = 32'o3524340615 ^ 32'o13402166523;
      8'b10010000: dzhxQnrxzS = 32'o11236155035 ^ 32'd293646697 ^ 32'o3250243652;
      8'hec: dzhxQnrxzS = 32'b00110010010011001011111111010100 ^ 32'd1930793738;
      8'b00100011: dzhxQnrxzS = 32'd3327297106 ^ 32'h872baa8c;
      8'd240: dzhxQnrxzS = 32'o23701257014 ^ 32'b11011110010111000111001011010010;
      8'd183: dzhxQnrxzS = 32'd2786597163 ^ 32'd2210736984 ^ 32'o14441017255;
      8'o71: dzhxQnrxzS = 32'h2ff2182c ^ 32'h6e8b34f2;
      8'o33: dzhxQnrxzS = 32'b01010110100110101101001001011111 ^ 32'd398720641;
      8'o153: dzhxQnrxzS = 32'd1199543464 ^ 32'b00000110001001101011100001110110;
      8'h7c: dzhxQnrxzS = 32'b11011111010110100100101101101100 ^ 32'b10011110000000110110011110110010;
      8'b00101101: dzhxQnrxzS = 32'h18254c45 ^ 32'hf3f8dfd6 ^ 32'd2862923597;
      8'o236: dzhxQnrxzS = 32'h74094b41 ^ 32'b00110101010100000110011110011111;
      8'o162: dzhxQnrxzS = 32'o27031544302 ^ 32'o37117762034;
      8'b01010100: dzhxQnrxzS = 32'b10100101110001001101100001000010 ^ 32'd3835557020;
      8'b10101010: dzhxQnrxzS = 32'd390423964 ^ 32'o12617044502;
      8'd212: dzhxQnrxzS = 32'd2001011044 ^ 32'he06a5809 ^ 32'b11010110011101100111010110110011;
      8'o105: dzhxQnrxzS = 32'b10111101100111100001000110010000 ^ 32'hfcc73d4e;
      8'o310: dzhxQnrxzS = 32'o34352215506 ^ 32'ha2f03798;
      8'd113: dzhxQnrxzS = 32'd664213186 ^ 32'd3897295006 ^ 32'o21640435202;
      8'b01110111: dzhxQnrxzS = 32'd2082671891 ^ 32'o37323311536 ^ 32'b11000110001101111011001010010011;
      8'hd0: dzhxQnrxzS = 32'd4002317018 ^ 32'b10111110010001010000000010111001 ^ 32'h1192aebd;
      8'o213: dzhxQnrxzS = 32'd4249495106 ^ 32'b10111100001100110000101010011100;
      8'o130: dzhxQnrxzS = 32'o20237104306 ^ 32'h50b05855 ^ 32'o22345376115;
      8'h7a: dzhxQnrxzS = 32'hfca6fb3 ^ 32'h483c1757 ^ 32'o653652072;
      8'ha1: dzhxQnrxzS = 32'hcd005140 ^ 32'd2356772254;
      8'd82: dzhxQnrxzS = 32'o11743323110 ^ 32'o1665105226;
      8'o233: dzhxQnrxzS = 32'o10200674710 ^ 32'o3031403425 ^ 32'h1b3c5203;
      8'd86: dzhxQnrxzS = 32'ha15b96d ^ 32'o11323112663;
      8'o31: dzhxQnrxzS = 32'o31156200240 ^ 32'h88c02c7e;
      8'hfb: dzhxQnrxzS = 32'd1712311847 ^ 32'd2603855251 ^ 32'b10111100011001010100111101101010;
      8'd219: dzhxQnrxzS = 32'd3692259940 ^ 32'b10011101010010100100011010111010;
      8'b11000111: dzhxQnrxzS = 32'he8020518 ^ 32'd2155214886 ^ 32'o5113550740;
      8'ha: dzhxQnrxzS = 32'd3648167983 ^ 32'o23002706361;
      8'h92: dzhxQnrxzS = 32'd2713734544 ^ 32'd4237793811 ^ 32'b00011100000011101111101101011101;
      8'hca: dzhxQnrxzS = 32'o14707441011 ^ 32'o3236235404 ^ 32'h3c3e55d3;
      8'o15: dzhxQnrxzS = 32'o12776650102 ^ 32'o2640476234;
      8'b01011010: dzhxQnrxzS = 32'd1297169986 ^ 32'd201855644;
      8'b10101101: dzhxQnrxzS = 32'o740165622 ^ 32'o20526676445 ^ 32'hc3a2ba69;
      8'd73: dzhxQnrxzS = 32'd3486694496 ^ 32'o21642710276;
      8'd48: dzhxQnrxzS = 32'b01000111000000011111011001000011 ^ 32'b00000110010110001101101010011101;
      8'o45: dzhxQnrxzS = 32'o4041073422 ^ 32'd1643994060;
      8'h70: dzhxQnrxzS = 32'o27503431546 ^ 32'hfc571fb8;
      8'hcc: dzhxQnrxzS = 32'o32556030360 ^ 32'b10010100111000010001110000101110;
      8'h8: dzhxQnrxzS = 32'hb1cdc9ad ^ 32'd4038387059;
      8'o42: dzhxQnrxzS = 32'hd0606397 ^ 32'd2436452169;
      8'h9f: dzhxQnrxzS = 32'd3745353052 ^ 32'h18338aa9 ^ 32'd2253859627;
      8'h5d: dzhxQnrxzS = 32'h72281d2f ^ 32'd863056369;
      8'b00000001: dzhxQnrxzS = 32'd3055059698 ^ 32'o4552125201 ^ 32'o32262202255;
      8'b10111000: dzhxQnrxzS = 32'd311448656 ^ 32'd1407809678;
      8'o140: dzhxQnrxzS = 32'o26672506023 ^ 32'b11001110110000000001000010110000 ^ 32'h3973b07d;
      8'b10000111: dzhxQnrxzS = 32'b11010101110110101100001001001001 ^ 32'b10010100101000111110111010010111;
      8'o200: dzhxQnrxzS = 32'o34163210244 ^ 32'b10111001111011110111110001111110 ^ 32'b00011001011110110100000000000100;
      8'b10101011: dzhxQnrxzS = 32'b01010100001111110000001011101100 ^ 32'd58202684 ^ 32'o2617432016;
      8'o115: dzhxQnrxzS = 32'b00010001011010000100000010100110 ^ 32'o5255624704 ^ 32'h7a8645bc;
      8'o46: dzhxQnrxzS = 32'o13530070776 ^ 32'o3416256440;
      8'b10000110: dzhxQnrxzS = 32'hf04e928 ^ 32'b01001110010111011100010111110110;
      8'd194: dzhxQnrxzS = 32'ha531c12b ^ 32'o26636767447 ^ 32'o12204601322;
      8'b10001111: dzhxQnrxzS = 32'b11110011011001111000100101110000 ^ 32'hb21ea5ae;
      8'hee: dzhxQnrxzS = 32'hfaef1884 ^ 32'b11010010111010111011101100101001 ^ 32'b01101001010111011000111101110011;
      8'd188: dzhxQnrxzS = 32'o5232717066 ^ 32'd1798484712;
      8'o344: dzhxQnrxzS = 32'b00010101010111111100100010100101 ^ 32'd1409737851;
      8'hc6: dzhxQnrxzS = 32'd4062273371 ^ 32'o26336071605;
      8'b00110101: dzhxQnrxzS = 32'o5342757 ^ 32'b00110100101000011100110101010010 ^ 32'd1976378467;
      8'b00011000: dzhxQnrxzS = 32'd4266358538 ^ 32'd990698331 ^ 32'b10000100001111101000000010001111;
      8'd222: dzhxQnrxzS = 32'd583933793 ^ 32'h44409963 ^ 32'o4765725334;
      8'b10110110: dzhxQnrxzS = 32'o35304357604 ^ 32'o25222171532;
    endcase
  end

  always_ff @(posedge clk_i) begin
    if(rst_i) begin
      Vx0I4zbHz <= '0;
    end
    else if (cSJpl8RGMw2bgs48nEfg[32'o11350642577 ^ 32'h4ba3456d]) begin
      Vx0I4zbHz <= '0;
    end
    else if(dNVOskLQGaCf26HqGY[32'd4176352419 ^ 32'o37073412241]) begin
      case(Pn7J)
        32'h00: Vx0I4zbHz <= data;
        32'h04: Vx0I4zbHz <= valid;
        32'h08: Vx0I4zbHz <= busy;
        32'h0c: Vx0I4zbHz <= baudrate;
        32'h10: Vx0I4zbHz <= parity_en;
        32'h14: Vx0I4zbHz <= stopbit;
        default: Vx0I4zbHz <= Vx0I4zbHz;
      endcase
    end
    else begin
      Vx0I4zbHz <= Vx0I4zbHz;
    end
  end

  always_ff @(posedge clk_i) begin
    if(rst_i) begin
      valid <= '0;
    end
    else begin
      valid <= dzhxQnrxzS[32'h281afbe5 ^ 32'd672857072];
    end
  end

  always_comb begin
    case ({CLD6rGMxYQM8yZ4, HWEbwjZ7R, raRSSx568gLgRd, C8sfwwEjm50H, N6jQMBhCLQ, sTe2Bcb7nHzYdOot, LhC})
      7'h68: yqfsQ7Rv18I3yx8 = 32'o30455604317 ^ 32'd2354701017 ^ 32'o17621670;
      7'o52: yqfsQ7Rv18I3yx8 = 32'b10100110001010111010100011011010 ^ 32'b10001011011110001111000101101110 ^ 32'h6582901a;
      7'o1: yqfsQ7Rv18I3yx8 = 32'o25035546667 ^ 32'd283310341 ^ 32'b11110000010001011111110100011100;
      7'b0010101: yqfsQ7Rv18I3yx8 = 32'o35022321533 ^ 32'o11731455103 ^ 32'b11101111111111100011000010110110;
      7'd56: yqfsQ7Rv18I3yx8 = 32'd3462099929 ^ 32'b10000110100010101011101001110111;
      7'd55: yqfsQ7Rv18I3yx8 = 32'd371011243 ^ 32'o36103510630 ^ 32'hafc2769d;
      7'h52: yqfsQ7Rv18I3yx8 = 32'd3992744870 ^ 32'hdf26d0a9 ^ 32'b01111010000010110110101010100001;
      7'o63: yqfsQ7Rv18I3yx8 = 32'b01101101110010010111011110101001 ^ 32'hd8021eeb ^ 32'o37506520354;
      7'b0001000: yqfsQ7Rv18I3yx8 = 32'b01001011001101110010101101011000 ^ 32'd137575865 ^ 32'd198565711;
      7'h21: yqfsQ7Rv18I3yx8 = 32'b01001100101111000010100011001011 ^ 32'd74309989;
      7'o113: yqfsQ7Rv18I3yx8 = 32'b00101101101011000011111010010011 ^ 32'o33526034340 ^ 32'b10111000001001011100111111011101;
      7'd34: yqfsQ7Rv18I3yx8 = 32'o20551477371 ^ 32'o31535733527;
      7'b0110010: yqfsQ7Rv18I3yx8 = 32'b10001001011011001100000010001010 ^ 32'd404175240 ^ 32'hd9aa30ac;
      7'o123: yqfsQ7Rv18I3yx8 = 32'o23552755037 ^ 32'd3581547441;
      7'o33: yqfsQ7Rv18I3yx8 = 32'b10001111010111000010111011100000 ^ 32'hbf629af ^ 32'd3430665953;
      7'h44: yqfsQ7Rv18I3yx8 = 32'b01010010000101101001100111100011 ^ 32'o3261650115;
      7'o171: yqfsQ7Rv18I3yx8 = 32'b10111011011011000100001001100100 ^ 32'o24635360433 ^ 32'h55c86ad0;
      7'h16: yqfsQ7Rv18I3yx8 = 32'd69600478 ^ 32'o31027146113 ^ 32'b10000100101010110000000100111011;
      7'h13: yqfsQ7Rv18I3yx8 = 32'b01111111111000010001110110000110 ^ 32'h3730d428;
      7'b1111110: yqfsQ7Rv18I3yx8 = 32'd1784541974 ^ 32'b11011011010111011001011111100100 ^ 32'd4191268188;
      7'o53: yqfsQ7Rv18I3yx8 = 32'o17157332260 ^ 32'hb56962ed ^ 32'b10000100000001010001111111110011;
      7'hb: yqfsQ7Rv18I3yx8 = 32'o33006662401 ^ 32'b10010000110010101010110010101111;
      7'b0101110: yqfsQ7Rv18I3yx8 = 32'o21043443346 ^ 32'd1540036149 ^ 32'h9b94997d;
      7'o124: yqfsQ7Rv18I3yx8 = 32'hd5edabaa ^ 32'h1f8ebedb ^ 32'd2192760031;
      7'd13: yqfsQ7Rv18I3yx8 = 32'o17210220342 ^ 32'b00110010111100001110100101001100;
      7'h62: yqfsQ7Rv18I3yx8 = 32'b10100110100110101011100111011111 ^ 32'd294549310 ^ 32'o37761203517;
      7'h3b: yqfsQ7Rv18I3yx8 = 32'd1211670747 ^ 32'd15296885;
      7'b1100000: yqfsQ7Rv18I3yx8 = 32'd804968885 ^ 32'h672b101b;
      7'd31: yqfsQ7Rv18I3yx8 = 32'b11101100010100110111001010011000 ^ 32'o16372075321 ^ 32'd3614097895;
      7'h19: yqfsQ7Rv18I3yx8 = 32'd1358406816 ^ 32'ha846898b ^ 32'hb060e485;
      7'd4: yqfsQ7Rv18I3yx8 = 32'o31431132140 ^ 32'd3601644767 ^ 32'o12206340421;
      7'o36: yqfsQ7Rv18I3yx8 = 32'hb2de6d7d ^ 32'd4285401662 ^ 32'b00000101011000011010111011101101;
      7'd40: yqfsQ7Rv18I3yx8 = 32'h383982a4 ^ 32'o16072045412;
      7'd79: yqfsQ7Rv18I3yx8 = 32'd68950775 ^ 32'd1288557401;
      7'b1110111: yqfsQ7Rv18I3yx8 = 32'd2844462574 ^ 32'he15ac440;
      7'b1111000: yqfsQ7Rv18I3yx8 = 32'o24755011655 ^ 32'd4016429571;
      7'o151: yqfsQ7Rv18I3yx8 = 32'o7730276106 ^ 32'o16754132750;
      7'o111: yqfsQ7Rv18I3yx8 = 32'b00100111001110011100000010101100 ^ 32'h6fe80902;
      7'o135: yqfsQ7Rv18I3yx8 = 32'h9b2a20b1 ^ 32'o5107557746 ^ 32'd4209325816;
      7'o0: yqfsQ7Rv18I3yx8 = 32'b10101101110100110001011100110010 ^ 32'o5513011767 ^ 32'hc82ecd6b;
      7'b1001100: yqfsQ7Rv18I3yx8 = 32'd2294071177 ^ 32'd3228399143;
      7'b1000101: yqfsQ7Rv18I3yx8 = 32'h95889f1d ^ 32'd1508994571 ^ 32'd2225617080;
      7'd52: yqfsQ7Rv18I3yx8 = 32'o24327670606 ^ 32'b11101011100011101011100000101000;
      7'd15: yqfsQ7Rv18I3yx8 = 32'd546571524 ^ 32'b10101001001010000011101111011111 ^ 32'o30133373565;
      7'o46: yqfsQ7Rv18I3yx8 = 32'o24014577000 ^ 32'd3907205038;
      7'o2: yqfsQ7Rv18I3yx8 = 32'd82288056 ^ 32'd2673537141 ^ 32'b11010011011011001010010001100011;
      7'b1111010: yqfsQ7Rv18I3yx8 = 32'd3368051195 ^ 32'b10000000000100011010100001010101;
      7'o12: yqfsQ7Rv18I3yx8 = 32'd968796802 ^ 32'b11000001000101101011000100111001 ^ 32'b10110000011110011101001000010101;
      7'o155: yqfsQ7Rv18I3yx8 = 32'd1753668384 ^ 32'h2057128e;
      7'o132: yqfsQ7Rv18I3yx8 = 32'd4058689830 ^ 32'd1258143510 ^ 32'd4089890718;
      7'o112: yqfsQ7Rv18I3yx8 = 32'd201050993 ^ 32'd1126826719;
      7'd5: yqfsQ7Rv18I3yx8 = 32'o21515403751 ^ 32'o22560405160 ^ 32'b01010000001001011100010000110111;
      7'h5c: yqfsQ7Rv18I3yx8 = 32'hc979e332 ^ 32'd2175281820;
      7'b1111111: yqfsQ7Rv18I3yx8 = 32'd3780067088 ^ 32'b01100100111101001001101001101100 ^ 32'b11001101011010100110110011010011;
      7'b1111011: yqfsQ7Rv18I3yx8 = 32'b10011100100000000111110100111110 ^ 32'd3596502773 ^ 32'b00000010000011111111001001100100;
      7'o156: yqfsQ7Rv18I3yx8 = 32'd456774884 ^ 32'b11001111100101001010011100101100 ^ 32'd2625419878;
      7'd39: yqfsQ7Rv18I3yx8 = 32'b11101101111101011110001001101110 ^ 32'd2770611136;
      7'o120: yqfsQ7Rv18I3yx8 = 32'b11100011001011110101010011000001 ^ 32'd2885590383;
      7'o145: yqfsQ7Rv18I3yx8 = 32'o10070544124 ^ 32'b00001000001100110000000111111010;
      7'b0011000: yqfsQ7Rv18I3yx8 = 32'b01010000110100100000000100000000 ^ 32'b00011000000000111100100010101110;
      7'b0000011: yqfsQ7Rv18I3yx8 = 32'd2311313672 ^ 32'o17470261447 ^ 32'o27574671601;
      7'h23: yqfsQ7Rv18I3yx8 = 32'o11744244572 ^ 32'o720100324;
      7'b0001001: yqfsQ7Rv18I3yx8 = 32'hd687f64 ^ 32'b01000101101110011011011011001010;
      7'o125: yqfsQ7Rv18I3yx8 = 32'b11000111110111101011000110111010 ^ 32'h8f0f7814;
      7'd45: yqfsQ7Rv18I3yx8 = 32'd169828432 ^ 32'o10263524776;
      7'h74: yqfsQ7Rv18I3yx8 = 32'd439545817 ^ 32'd1390618231;
      7'b1001110: yqfsQ7Rv18I3yx8 = 32'd3297649394 ^ 32'b10001100010111111110101101011100;
      7'd37: yqfsQ7Rv18I3yx8 = 32'o33625624672 ^ 32'o20201630615 ^ 32'h1481d199;
      7'd49: yqfsQ7Rv18I3yx8 = 32'hedc2b908 ^ 32'o24504670246;
      7'h3f: yqfsQ7Rv18I3yx8 = 32'b01100110110110011001001110000100 ^ 32'o25121253552 ^ 32'd2269973824;
      7'b0111010: yqfsQ7Rv18I3yx8 = 32'b01011000100011110010011101111011 ^ 32'd274656981;
      7'h17: yqfsQ7Rv18I3yx8 = 32'd76643028 ^ 32'ha13eb1a7 ^ 32'o35537401335;
      7'o60: yqfsQ7Rv18I3yx8 = 32'd577737349 ^ 32'b01101010101111100101101100101011;
      7'h6c: yqfsQ7Rv18I3yx8 = 32'o12021564174 ^ 32'b00011000100101110010000111010010;
      7'd103: yqfsQ7Rv18I3yx8 = 32'b01100001110000100111001111011100 ^ 32'd689158770;
      7'd100: yqfsQ7Rv18I3yx8 = 32'b00010001001111001100011100010000 ^ 32'b01011001111011010000111010111110;
      7'h3c: yqfsQ7Rv18I3yx8 = 32'h982ab239 ^ 32'o6127156101 ^ 32'he1a7a7d6;
      7'o44: yqfsQ7Rv18I3yx8 = 32'd3972210945 ^ 32'd2752702639;
      7'd106: yqfsQ7Rv18I3yx8 = 32'd440202062 ^ 32'd667684803 ^ 32'd1965110563;
      7'd61: yqfsQ7Rv18I3yx8 = 32'd3506594592 ^ 32'h99d3aa8e;
      7'h71: yqfsQ7Rv18I3yx8 = 32'h4437bf33 ^ 32'd1746520354 ^ 32'h64ffbfbf;
      7'd107: yqfsQ7Rv18I3yx8 = 32'h540e1fc8 ^ 32'd484431462;
      7'd99: yqfsQ7Rv18I3yx8 = 32'heb926cf8 ^ 32'd2739119446;
      7'b1011110: yqfsQ7Rv18I3yx8 = 32'h9e191068 ^ 32'd3677931408 ^ 32'b00001101111100000001111001010110;
      7'h14: yqfsQ7Rv18I3yx8 = 32'h274e5401 ^ 32'o15747716657;
      7'h66: yqfsQ7Rv18I3yx8 = 32'b10010011101111001001100100100110 ^ 32'b10001001000110100010111111101110 ^ 32'd1383563110;
      7'o141: yqfsQ7Rv18I3yx8 = 32'd2847358924 ^ 32'b11010101000111011001101000010011 ^ 32'b00110100011110110110110001110001;
      7'h42: yqfsQ7Rv18I3yx8 = 32'o6104125535 ^ 32'h2293eca0 ^ 32'o13324507123;
      7'o100: yqfsQ7Rv18I3yx8 = 32'd1926214185 ^ 32'h3a1e7b87;
      7'h1c: yqfsQ7Rv18I3yx8 = 32'h5e6681e5 ^ 32'b00010110101101110100100001001011;
      7'h43: yqfsQ7Rv18I3yx8 = 32'o12524576362 ^ 32'd991812500 ^ 32'h269eeec8;
      7'b1011001: yqfsQ7Rv18I3yx8 = 32'b01010110101100000011111101000101 ^ 32'b00011110011000011111011011101010;
      7'b0000111: yqfsQ7Rv18I3yx8 = 32'o35601621123 ^ 32'b10100110110101101110101111111101;
      7'o20: yqfsQ7Rv18I3yx8 = 32'o27432021042 ^ 32'd4105825164;
      7'o165: yqfsQ7Rv18I3yx8 = 32'o26702315245 ^ 32'hffd8530b;
      7'd26: yqfsQ7Rv18I3yx8 = 32'd990619226 ^ 32'h5ade37a2 ^ 32'h29045856;
      7'o107: yqfsQ7Rv18I3yx8 = 32'd1881648976 ^ 32'd955672318;
      7'o57: yqfsQ7Rv18I3yx8 = 32'h2898d161 ^ 32'hce6603b2 ^ 32'o25613615575;
      7'o121: yqfsQ7Rv18I3yx8 = 32'd2922680297 ^ 32'h96f17b51 ^ 32'h70143d16;
      7'd57: yqfsQ7Rv18I3yx8 = 32'o24423521064 ^ 32'o20016106374 ^ 32'o15451763546;
      7'o51: yqfsQ7Rv18I3yx8 = 32'b11110000010100000111010010100101 ^ 32'd1967273439 ^ 32'b11001101110000111000100011010100;
      7'd70: yqfsQ7Rv18I3yx8 = 32'o35526511571 ^ 32'b10010111010100101001100111101110 ^ 32'd853132089;
      7'o160: yqfsQ7Rv18I3yx8 = 32'd3302181846 ^ 32'd2348974712;
      7'h12: yqfsQ7Rv18I3yx8 = 32'hf1842b69 ^ 32'b10111001010101011110001011000111;
      7'b0111110: yqfsQ7Rv18I3yx8 = 32'b10111110110011110001011100111000 ^ 32'b11110110000111101101111010010110;
      7'o133: yqfsQ7Rv18I3yx8 = 32'd4102955092 ^ 32'b10111100010111111110100111111011;
      7'h6: yqfsQ7Rv18I3yx8 = 32'b01100001100111100001111110010010 ^ 32'd693098044;
      7'd124: yqfsQ7Rv18I3yx8 = 32'he9076095 ^ 32'o24165524473;
      7'd32: yqfsQ7Rv18I3yx8 = 32'h741ade04 ^ 32'o7462613652;
      7'o157: yqfsQ7Rv18I3yx8 = 32'd1035421527 ^ 32'd1969655545;
      7'd72: yqfsQ7Rv18I3yx8 = 32'b10101000110100011100100010000100 ^ 32'd3758096682;
      7'd44: yqfsQ7Rv18I3yx8 = 32'b01100001101111010011000000010010 ^ 32'b11011100111111111001110000010001 ^ 32'd4120077741;
      7'd87: yqfsQ7Rv18I3yx8 = 32'o20417645167 ^ 32'hccee83d9;
      7'd115: yqfsQ7Rv18I3yx8 = 32'd1287566423 ^ 32'd74415609;
      7'b0001100: yqfsQ7Rv18I3yx8 = 32'o27062240203 ^ 32'd4028139821;
      7'b1001101: yqfsQ7Rv18I3yx8 = 32'o21337675464 ^ 32'b11100100111111010110011010110111 ^ 32'b00100111010100111101010000101101;
      7'h1d: yqfsQ7Rv18I3yx8 = 32'b11100010111101110010011000001000 ^ 32'd2854678438;
      7'h76: yqfsQ7Rv18I3yx8 = 32'hea72c0fd ^ 32'd1379131502 ^ 32'd4036028733;
      7'd114: yqfsQ7Rv18I3yx8 = 32'h5043032d ^ 32'b00011000100100101100101010000011;
      7'h56: yqfsQ7Rv18I3yx8 = 32'd2264426144 ^ 32'o31612327416;
      7'd53: yqfsQ7Rv18I3yx8 = 32'o13626764637 ^ 32'b00101111011000010101100010100011 ^ 32'h39eb7892;
      7'o137: yqfsQ7Rv18I3yx8 = 32'h6dbd1102 ^ 32'b01100101000000110111111100100000 ^ 32'b01000000011011111010011110001101;
      7'd125: yqfsQ7Rv18I3yx8 = 32'd2966557240 ^ 32'o21447743405 ^ 32'h749c1c92;
      7'd88: yqfsQ7Rv18I3yx8 = 32'b01001000001000011101111010000010 ^ 32'b00000000111100000001011100101100;
      7'd54: yqfsQ7Rv18I3yx8 = 32'd4145840102 ^ 32'd3217929800;
      7'o16: yqfsQ7Rv18I3yx8 = 32'd863013938 ^ 32'h14f42824 ^ 32'b01101111010101010110110110111000;
      7'o21: yqfsQ7Rv18I3yx8 = 32'o37653643370 ^ 32'd3260654023 ^ 32'd1948724881;
      7'b1000001: yqfsQ7Rv18I3yx8 = 32'hc9cc9154 ^ 32'b01100101011011111001101010010010 ^ 32'b11100100011100101100001001101000;
    endcase
  end

  logic [31:0] vKAzElEBQ5fg3z;
  always_comb begin
    case ({LhC, raRSSx568gLgRd, sTe2Bcb7nHzYdOot, CLD6rGMxYQM8yZ4, HWEbwjZ7R, N6jQMBhCLQ, C8sfwwEjm50H})
      7'b1111011: vKAzElEBQ5fg3z = 32'd80571196 ^ 32'd478445144 ^ 32'o17463462625;
      7'd94: vKAzElEBQ5fg3z = 32'h26651b5d ^ 32'b01000010111000100110101110101100;
      7'hb: vKAzElEBQ5fg3z = 32'd2665906835 ^ 32'hfa61f262;
      7'h79: vKAzElEBQ5fg3z = 32'o25701775556 ^ 32'h28eff04 ^ 32'he90e749b;
      7'b1100000: vKAzElEBQ5fg3z = 32'o1176355365 ^ 32'b10000001011011111111011101110011 ^ 32'hcc115d77;
      7'o54: vKAzElEBQ5fg3z = 32'd4254298845 ^ 32'o16033711204 ^ 32'hc97b90a8;
      7'h14: vKAzElEBQ5fg3z = 32'b11011010110001110001100101111110 ^ 32'h4e333d06 ^ 32'o32034652211;
      7'd105: vKAzElEBQ5fg3z = 32'o16266307334 ^ 32'b00111000100101110001000111111010 ^ 32'hec9efd7;
      7'h11: vKAzElEBQ5fg3z = 32'b10011001000011011011001001110010 ^ 32'd3716858499;
      7'd115: vKAzElEBQ5fg3z = 32'd2036471931 ^ 32'h1184ff87 ^ 32'd207722253;
      7'h3f: vKAzElEBQ5fg3z = 32'h172e2504 ^ 32'o16352252765;
      7'b0000110: vKAzElEBQ5fg3z = 32'o35546747663 ^ 32'b11010110011010111011000100010001 ^ 32'b01011111011101110000111001010011;
      7'd22: vKAzElEBQ5fg3z = 32'b00100000111001011010011100101110 ^ 32'b10010111011101111000100011011111 ^ 32'hd3155f00;
      7'o66: vKAzElEBQ5fg3z = 32'b10011011110110011111010111110110 ^ 32'd338824066 ^ 32'heb6c8e85;
      7'o4: vKAzElEBQ5fg3z = 32'hccdce4de ^ 32'o30636511001 ^ 32'd1310787118;
      7'b0000011: vKAzElEBQ5fg3z = 32'd2630803461 ^ 32'd1155236504 ^ 32'b10111100100100100001001001101100;
      7'd103: vKAzElEBQ5fg3z = 32'b11101010000100011100111001000010 ^ 32'b10011011100111000001101100100010 ^ 32'o2502522621;
      7'h23: vKAzElEBQ5fg3z = 32'b10011110110010101111100111001001 ^ 32'hfa4d8938;
      7'b1011000: vKAzElEBQ5fg3z = 32'b10111011101110101010101000110011 ^ 32'b11111111001111011101101011000010;
      7'o45: vKAzElEBQ5fg3z = 32'b10101001110111011010101010111010 ^ 32'b11101101010110101101101001001011;
      7'h7f: vKAzElEBQ5fg3z = 32'd63664573 ^ 32'b11110000001110001100111011100101 ^ 32'o22735147651;
      7'd74: vKAzElEBQ5fg3z = 32'b11110001011010000100100101111001 ^ 32'o5104046537 ^ 32'd3170858199;
      7'o141: vKAzElEBQ5fg3z = 32'd3814128591 ^ 32'o24764305476;
      7'h17: vKAzElEBQ5fg3z = 32'b10110111110010100011010000010001 ^ 32'd1499594336 ^ 32'o21213135200;
      7'd107: vKAzElEBQ5fg3z = 32'b00010110010101010010010000010001 ^ 32'h51da3d75 ^ 32'o4302064625;
      7'h1a: vKAzElEBQ5fg3z = 32'o20672146662 ^ 32'b11000010110110001010010111110101 ^ 32'd548870326;
      7'b1111110: vKAzElEBQ5fg3z = 32'd4122659067 ^ 32'd3091679369 ^ 32'd695922819;
      7'o25: vKAzElEBQ5fg3z = 32'h33e54843 ^ 32'h776238b2;
      7'b0110001: vKAzElEBQ5fg3z = 32'h7c4016bd ^ 32'b00111000110001110110011001001100;
      7'b0100100: vKAzElEBQ5fg3z = 32'b10001011100111111001011110011101 ^ 32'd3587931697 ^ 32'd449026397;
      7'b0110100: vKAzElEBQ5fg3z = 32'h3e175337 ^ 32'd2056266694;
      7'b1001011: vKAzElEBQ5fg3z = 32'd1456356993 ^ 32'hdaac2501 ^ 32'd3907349361;
      7'd33: vKAzElEBQ5fg3z = 32'd1447812703 ^ 32'h12ccaeae;
      7'b1000110: vKAzElEBQ5fg3z = 32'd302014487 ^ 32'd1988563174;
      7'd9: vKAzElEBQ5fg3z = 32'o25756665176 ^ 32'd1060915148 ^ 32'o32400056503;
      7'b1100110: vKAzElEBQ5fg3z = 32'o31716277315 ^ 32'b00110110101000100111001101010110 ^ 32'h9d1c7d6a;
      7'b0001010: vKAzElEBQ5fg3z = 32'b01000100000011010100001000110110 ^ 32'h208a32c7;
      7'h7c: vKAzElEBQ5fg3z = 32'd1040051221 ^ 32'b01010111100010111100010001001100 ^ 32'd787568808;
      7'd0: vKAzElEBQ5fg3z = 32'hc13db314 ^ 32'b01110110110111100011011010110101 ^ 32'b11110011011001001111010101010000;
      7'b0111101: vKAzElEBQ5fg3z = 32'd1446521610 ^ 32'd314530811;
      7'd16: vKAzElEBQ5fg3z = 32'h850ff1eb ^ 32'd559107191 ^ 32'o34066746555;
      7'b0100010: vKAzElEBQ5fg3z = 32'hf5e99f44 ^ 32'd3531631396 ^ 32'b01000011111011101000010010010001;
      7'o5: vKAzElEBQ5fg3z = 32'o15521170274 ^ 32'h29c3804d;
      7'h7d: vKAzElEBQ5fg3z = 32'ha0517359 ^ 32'he4d603a8;
      7'o155: vKAzElEBQ5fg3z = 32'o4154245677 ^ 32'hea7246cc ^ 32'h8f447d82;
      7'o165: vKAzElEBQ5fg3z = 32'b01110001000010110111001100010011 ^ 32'o12447225413 ^ 32'd1628514537;
      7'b0011000: vKAzElEBQ5fg3z = 32'h3607faab ^ 32'd2200026261 ^ 32'hf1a136cf;
      7'o55: vKAzElEBQ5fg3z = 32'o36136346220 ^ 32'b10110101111111101011110001100001;
      7'o117: vKAzElEBQ5fg3z = 32'b11011011011111000001000101111101 ^ 32'b10011011110000011101101010101001 ^ 32'o4416535445;
      7'h5b: vKAzElEBQ5fg3z = 32'o7125525515 ^ 32'o656115006 ^ 32'd1533624762;
      7'b0101011: vKAzElEBQ5fg3z = 32'd1111651829 ^ 32'd650446084;
      7'b0100110: vKAzElEBQ5fg3z = 32'h49431f6b ^ 32'heae13e2b ^ 32'hc72551b1;
      7'h2e: vKAzElEBQ5fg3z = 32'o4377304624 ^ 32'o10736574545;
      7'd7: vKAzElEBQ5fg3z = 32'b00010000110111111101101110011101 ^ 32'o16722115673 ^ 32'o304030327;
      7'd56: vKAzElEBQ5fg3z = 32'd3952789935 ^ 32'o25707334536;
      7'b1001110: vKAzElEBQ5fg3z = 32'b00111110001000111100001111111000 ^ 32'b01011010101001001011001100001001;
      7'd71: vKAzElEBQ5fg3z = 32'hb2a0d693 ^ 32'd3719835716 ^ 32'd195008038;
      7'b0001111: vKAzElEBQ5fg3z = 32'o16037417272 ^ 32'd388964078 ^ 32'b00000011110101100111000010100101;
      7'b0111110: vKAzElEBQ5fg3z = 32'o3337716070 ^ 32'hbff83533 ^ 32'o30000154772;
      7'b1110001: vKAzElEBQ5fg3z = 32'had002fd3 ^ 32'h9a0b225e ^ 32'd1938587004;
      7'b0011100: vKAzElEBQ5fg3z = 32'o7464027447 ^ 32'h78575fd6;
      7'o114: vKAzElEBQ5fg3z = 32'd3654239622 ^ 32'b10011101010010000011010101110111;
      7'b0111100: vKAzElEBQ5fg3z = 32'h445c5df4 ^ 32'o30103607125 ^ 32'd3251905360;
      7'd2: vKAzElEBQ5fg3z = 32'o22715217716 ^ 32'b11110011101100100110111100111111;
      7'o23: vKAzElEBQ5fg3z = 32'd2143779749 ^ 32'd2199210336 ^ 32'b10011000010101010100001000110100;
      7'b0110000: vKAzElEBQ5fg3z = 32'heec57a1e ^ 32'd2856454895;
      7'o123: vKAzElEBQ5fg3z = 32'd1627621477 ^ 32'o4162023202 ^ 32'o4423157026;
      7'd101: vKAzElEBQ5fg3z = 32'b00001010110010100100001010110010 ^ 32'd1207025005 ^ 32'd163352366;
      7'o144: vKAzElEBQ5fg3z = 32'o10577251561 ^ 32'o35224642752 ^ 32'heb29666a;
      7'o15: vKAzElEBQ5fg3z = 32'o30723743705 ^ 32'd586346820 ^ 32'ha13a4670;
      7'h68: vKAzElEBQ5fg3z = 32'd1669763610 ^ 32'o4700361353;
      7'd31: vKAzElEBQ5fg3z = 32'b10100001100011111001011101011100 ^ 32'b11011100001001011100001110111001 ^ 32'o3113222024;
      7'b1011101: vKAzElEBQ5fg3z = 32'o15326050675 ^ 32'd2225362333 ^ 32'b10101011011110110111010011010001;
      7'h27: vKAzElEBQ5fg3z = 32'b11001001110111101011011101101010 ^ 32'd2531902076 ^ 32'b00111011101100000000010111100111;
      7'o16: vKAzElEBQ5fg3z = 32'h6af1a3e6 ^ 32'd242668311;
      7'h5f: vKAzElEBQ5fg3z = 32'b00100000111010011001010010000100 ^ 32'd1087912119 ^ 32'o455556302;
      7'h42: vKAzElEBQ5fg3z = 32'd84374112 ^ 32'h61800291;
      7'o121: vKAzElEBQ5fg3z = 32'h52136cd4 ^ 32'o2645016045;
      7'h7a: vKAzElEBQ5fg3z = 32'o23215616304 ^ 32'hfeb06c35;
      7'h54: vKAzElEBQ5fg3z = 32'd185316470 ^ 32'b10001011011101101010010110111001 ^ 32'd3304743230;
      7'b1110111: vKAzElEBQ5fg3z = 32'b11110110101001111110010011101110 ^ 32'b10010010001000001001010000011111;
      7'h5a: vKAzElEBQ5fg3z = 32'd3088546922 ^ 32'hdc900c9b;
      7'd67: vKAzElEBQ5fg3z = 32'd2343575266 ^ 32'o5343557642 ^ 32'hc4b9b1b1;
      7'b0111011: vKAzElEBQ5fg3z = 32'o26540166463 ^ 32'o32101716702;
      7'h78: vKAzElEBQ5fg3z = 32'd2006700077 ^ 32'd3456731005 ^ 32'd4246022049;
      7'h4d: vKAzElEBQ5fg3z = 32'd2288811888 ^ 32'hcceb0f81;
      7'h76: vKAzElEBQ5fg3z = 32'h2ec8391e ^ 32'o20266247177 ^ 32'hc8960790;
      7'h19: vKAzElEBQ5fg3z = 32'o4017452662 ^ 32'hf311bb3c ^ 32'd2544410239;
      7'h33: vKAzElEBQ5fg3z = 32'b11100010111101011001110000010010 ^ 32'd2505472984 ^ 32'h1324973b;
      7'o122: vKAzElEBQ5fg3z = 32'h3d588c1b ^ 32'd925677324 ^ 32'd1861438438;
      7'd27: vKAzElEBQ5fg3z = 32'h7b4651a2 ^ 32'b10101111110101000011101011110000 ^ 32'o26005215643;
      7'd1: vKAzElEBQ5fg3z = 32'h60124713 ^ 32'b00100100100101010011011111100010;
      7'b0110010: vKAzElEBQ5fg3z = 32'h58f18f0b ^ 32'h3c76fffa;
      7'b0011101: vKAzElEBQ5fg3z = 32'hbbac1fdf ^ 32'o15133161436 ^ 32'o22621706060;
      7'o105: vKAzElEBQ5fg3z = 32'he2281a36 ^ 32'd2796513991;
      7'd99: vKAzElEBQ5fg3z = 32'b10111100000011011111011001101010 ^ 32'b01110100001101100010100110011101 ^ 32'b10101100101111001010111100000110;
      7'o164: vKAzElEBQ5fg3z = 32'b11011011110010111010100100111110 ^ 32'd1905931880 ^ 32'b11101110110101101110111110100111;
      7'b1010101: vKAzElEBQ5fg3z = 32'b00110101101010110001001001101001 ^ 32'o27346512615 ^ 32'hcab6f715;
      7'o100: vKAzElEBQ5fg3z = 32'b11001011011010011000111100000001 ^ 32'o21773577760;
      7'h29: vKAzElEBQ5fg3z = 32'o22046406160 ^ 32'b10011011011000011100010011110100 ^ 32'h4f7cb875;
      7'h2a: vKAzElEBQ5fg3z = 32'b00001101001000011110101000101110 ^ 32'h3fece6f4 ^ 32'b01010110010010100111110000101011;
      7'd40: vKAzElEBQ5fg3z = 32'o23133475702 ^ 32'b00100011101011011011110110011101 ^ 32'o37621133256;
      7'hc: vKAzElEBQ5fg3z = 32'b10101011000110011000111011011011 ^ 32'b11101111100111101111111000101010;
      7'h3a: vKAzElEBQ5fg3z = 32'o35025635534 ^ 32'b10001100110100000100101110101101;
      7'h1e: vKAzElEBQ5fg3z = 32'o27670350131 ^ 32'o33231520250;
      7'h6e: vKAzElEBQ5fg3z = 32'd806505637 ^ 32'b11000101111011000001010011110101 ^ 32'h917928a1;
      7'd65: vKAzElEBQ5fg3z = 32'hb7056418 ^ 32'o12123425426 ^ 32'b10100010110011000011111111111111;
      7'd114: vKAzElEBQ5fg3z = 32'd352601357 ^ 32'b01110001100000110011010111111100;
      7'd112: vKAzElEBQ5fg3z = 32'o13271575216 ^ 32'h1e618a7f;
      7'o131: vKAzElEBQ5fg3z = 32'o22271465001 ^ 32'o32630215360;
      7'd32: vKAzElEBQ5fg3z = 32'o31614546032 ^ 32'h84f56e19 ^ 32'o1620151362;
      7'd98: vKAzElEBQ5fg3z = 32'd575952546 ^ 32'b01111011100010101001100010000111 ^ 32'h3d59bed4;
      7'h6f: vKAzElEBQ5fg3z = 32'o6667522513 ^ 32'h5259d5ba;
      7'h8: vKAzElEBQ5fg3z = 32'h87a0cc85 ^ 32'o30356341301 ^ 32'd10387125;
      7'o65: vKAzElEBQ5fg3z = 32'd2835900992 ^ 32'o6042135344 ^ 32'd3708264533;
      7'b1010111: vKAzElEBQ5fg3z = 32'd3048519375 ^ 32'd3509831230;
      7'b0010010: vKAzElEBQ5fg3z = 32'd2473485214 ^ 32'o36772211557;
      7'b1010000: vKAzElEBQ5fg3z = 32'd4252754047 ^ 32'hf9261885 ^ 32'b01000000110110101000100000001011;
      7'h48: vKAzElEBQ5fg3z = 32'b11110001000101110001001101001101 ^ 32'd3282912822 ^ 32'h763d258a;
      7'b1010110: vKAzElEBQ5fg3z = 32'o33742762077 ^ 32'hbb0c94ce;
      7'b1001001: vKAzElEBQ5fg3z = 32'b01111111100000110110011111100110 ^ 32'h3b041717;
      7'h37: vKAzElEBQ5fg3z = 32'b11101010111101101000110100101001 ^ 32'b11110011000111000011000100000110 ^ 32'd2104347870;
      7'd106: vKAzElEBQ5fg3z = 32'd23405832 ^ 32'h6a85fb6d ^ 32'hf67ae94;
      7'h6c: vKAzElEBQ5fg3z = 32'hb93ed413 ^ 32'h716e8759 ^ 32'h8cd723bb;
      7'b0101111: vKAzElEBQ5fg3z = 32'hedb5f2b4 ^ 32'o1404754063 ^ 32'h85215a76;
      7'd57: vKAzElEBQ5fg3z = 32'd997927310 ^ 32'o17777054577;
      7'o104: vKAzElEBQ5fg3z = 32'h547990e5 ^ 32'o2077560024;
      7'b1011100: vKAzElEBQ5fg3z = 32'd1971331364 ^ 32'b00110001000001110101000111010101;
    endcase
  end

  assign CLD6rGMxYQM8yZ4 = Pn7J == (32'h325bfce8 ^ 32'b01000000011000001010001001001010 ^ 32'd1916493446);
  always_ff @(posedge clk_i) begin
    if(rst_i) begin
      data <= '0;
    end else if (yqfsQ7Rv18I3yx8[32'd3000100153 ^ 32'b10110010110100011110010100111001]) begin
      data <= '0;
    end
    else if(vKAzElEBQ5fg3z[32'he3e71f6d ^ 32'b00010001010110100000101100000110 ^ 32'hf2bd1476]) begin
      data <= t26Xa3D9y;
    end
    else begin
      data <= data;
    end
  end

  logic jV8bIfqHdflwW;
  logic [31:0] w6aL01ok1NWMnhRdDAP;
  always_comb begin
    case ({LhC, raRSSx568gLgRd, CLD6rGMxYQM8yZ4, busy, jV8bIfqHdflwW, C8sfwwEjm50H})
      6'b101001: w6aL01ok1NWMnhRdDAP = 32'b00110111011111010100011111100111 ^ 32'h3127073a;
      6'o46: w6aL01ok1NWMnhRdDAP = 32'd502897647 ^ 32'h1ba3db32;
      6'o31: w6aL01ok1NWMnhRdDAP = 32'o31653300021 ^ 32'o23065402000 ^ 32'o12010342314;
      6'h6: w6aL01ok1NWMnhRdDAP = 32'b11010001110101100001110101100011 ^ 32'hd78c5dbe;
      6'o16: w6aL01ok1NWMnhRdDAP = 32'h9ec6838c ^ 32'o23047141521;
      6'h1a: w6aL01ok1NWMnhRdDAP = 32'o24367755336 ^ 32'ha5859a03;
      6'd18: w6aL01ok1NWMnhRdDAP = 32'h82d12673 ^ 32'h82ff4dc7 ^ 32'o635025551;
      6'h36: w6aL01ok1NWMnhRdDAP = 32'o24736710214 ^ 32'b00000111000111100010111001100001 ^ 32'd2789211696;
      6'd5: w6aL01ok1NWMnhRdDAP = 32'b01001001111011011110101001100111 ^ 32'd937973129 ^ 32'd2019557171;
      6'o53: w6aL01ok1NWMnhRdDAP = 32'hcf1d03c9 ^ 32'hc9474314;
      6'h35: w6aL01ok1NWMnhRdDAP = 32'b01001010011101000111010001100111 ^ 32'b11001111011101110000101100101000 ^ 32'b10000011010110010011111110010010;
      6'h1: w6aL01ok1NWMnhRdDAP = 32'd1166904454 ^ 32'o10365746133;
      6'd57: w6aL01ok1NWMnhRdDAP = 32'o30152424547 ^ 32'o30774264672;
      6'd0: w6aL01ok1NWMnhRdDAP = 32'o22604665445 ^ 32'h90492bf8;
      6'o15: w6aL01ok1NWMnhRdDAP = 32'h7314d351 ^ 32'b11101010100011101011011111111010 ^ 32'b10011111110000000010010001110110;
      6'h24: w6aL01ok1NWMnhRdDAP = 32'o24222723417 ^ 32'o13707337444 ^ 32'd4211890422;
      6'o4: w6aL01ok1NWMnhRdDAP = 32'b00101111111011011001001101100010 ^ 32'o5155751677;
      6'd40: w6aL01ok1NWMnhRdDAP = 32'b11001000100110111110001110101001 ^ 32'd924113319 ^ 32'd4191517395;
      6'b111110: w6aL01ok1NWMnhRdDAP = 32'h71f45e1c ^ 32'h77ae1ec1;
      6'b100111: w6aL01ok1NWMnhRdDAP = 32'b11110000010000111101101100000100 ^ 32'b00100010011011010011101111100110 ^ 32'd3564412991;
      6'o45: w6aL01ok1NWMnhRdDAP = 32'hc61711c5 ^ 32'h31e84f1 ^ 32'o30324752751;
      6'd19: w6aL01ok1NWMnhRdDAP = 32'b00001010001111111010000011010111 ^ 32'o1431360012;
      6'b011100: w6aL01ok1NWMnhRdDAP = 32'b00101000110110101010110100110110 ^ 32'hc2780698 ^ 32'b11101100111110001110101101110011;
      6'h31: w6aL01ok1NWMnhRdDAP = 32'o32263617745 ^ 32'h6f294140 ^ 32'hbbbc1e78;
      6'h23: w6aL01ok1NWMnhRdDAP = 32'b11111000001101001101001010110100 ^ 32'hc1ac4145 ^ 32'd1069732652;
      6'd46: w6aL01ok1NWMnhRdDAP = 32'd1488437019 ^ 32'h5eedffc6;
      6'd30: w6aL01ok1NWMnhRdDAP = 32'd1486378396 ^ 32'o13660412501;
      6'd21: w6aL01ok1NWMnhRdDAP = 32'b00110100010100011110101011111010 ^ 32'b00110010000010111010101000100111;
      6'b010000: w6aL01ok1NWMnhRdDAP = 32'b11101101110001011110110101001011 ^ 32'b11101011100111111010110110010110;
      6'o60: w6aL01ok1NWMnhRdDAP = 32'o11772734157 ^ 32'o33164747734 ^ 32'o22030433556;
      6'o42: w6aL01ok1NWMnhRdDAP = 32'b01100001110001011000110110000010 ^ 32'd1368030168 ^ 32'h3615b687;
      6'o54: w6aL01ok1NWMnhRdDAP = 32'hab54868 ^ 32'd216991925;
      6'o13: w6aL01ok1NWMnhRdDAP = 32'o5153121532 ^ 32'b00101111111101101110001110000111;
      6'd32: w6aL01ok1NWMnhRdDAP = 32'h666706a7 ^ 32'o14017243172;
      6'b001100: w6aL01ok1NWMnhRdDAP = 32'ha77ae1b6 ^ 32'b10100001001000001010000101101011;
      6'b001001: w6aL01ok1NWMnhRdDAP = 32'b10111110001010101101111110100101 ^ 32'hb8709f78;
      6'h16: w6aL01ok1NWMnhRdDAP = 32'd1695615842 ^ 32'o14322645677;
      6'b110111: w6aL01ok1NWMnhRdDAP = 32'd4055162984 ^ 32'd791155832 ^ 32'o33061532315;
      6'hf: w6aL01ok1NWMnhRdDAP = 32'hc8075810 ^ 32'd3462207693;
      6'd56: w6aL01ok1NWMnhRdDAP = 32'o7002277352 ^ 32'd1045642807;
      6'h14: w6aL01ok1NWMnhRdDAP = 32'o5107147367 ^ 32'o27255612355 ^ 32'b10010101111100011001101011000111;
      6'b011101: w6aL01ok1NWMnhRdDAP = 32'hd3460df7 ^ 32'hd51c4d2a;
      6'b010111: w6aL01ok1NWMnhRdDAP = 32'd2369733286 ^ 32'b01010101001000000111100101100110 ^ 32'hde457b1d;
      6'h2a: w6aL01ok1NWMnhRdDAP = 32'd3081067190 ^ 32'b10110001111111110001101001101011;
      6'ha: w6aL01ok1NWMnhRdDAP = 32'o25160022321 ^ 32'h20d45c3c ^ 32'd2404268080;
      6'd60: w6aL01ok1NWMnhRdDAP = 32'hcd3e3893 ^ 32'd3063987814 ^ 32'b01111101110001001100011000101000;
      6'h3: w6aL01ok1NWMnhRdDAP = 32'h283462ba ^ 32'd778969703;
      6'd52: w6aL01ok1NWMnhRdDAP = 32'd1940981520 ^ 32'o16572643715;
      6'h1b: w6aL01ok1NWMnhRdDAP = 32'o26414500573 ^ 32'd1330724521 ^ 32'hfd39ff0f;
      6'o41: w6aL01ok1NWMnhRdDAP = 32'o35465106310 ^ 32'o642613072 ^ 32'o35401355057;
      6'b101101: w6aL01ok1NWMnhRdDAP = 32'hd0d3436f ^ 32'o15506301715 ^ 32'hbb90807f;
      6'h3a: w6aL01ok1NWMnhRdDAP = 32'o31203136277 ^ 32'b11001100010101101111110001100010;
      6'o77: w6aL01ok1NWMnhRdDAP = 32'hc3f7223 ^ 32'b00001010011001000011001011111110;
      6'h32: w6aL01ok1NWMnhRdDAP = 32'd1312786605 ^ 32'o11031344160;
      6'h3b: w6aL01ok1NWMnhRdDAP = 32'o26270144011 ^ 32'd3032189140;
      6'd61: w6aL01ok1NWMnhRdDAP = 32'o112137236 ^ 32'b11011010111101101110000101001011 ^ 32'hdd851f08;
      6'o57: w6aL01ok1NWMnhRdDAP = 32'o6325173665 ^ 32'h484d26b7 ^ 32'o17520710737;
      6'b011000: w6aL01ok1NWMnhRdDAP = 32'o22520072576 ^ 32'o5253112255 ^ 32'd3115753742;
      6'd8: w6aL01ok1NWMnhRdDAP = 32'hdfbb4323 ^ 32'b11011001111000010000001111111110;
      6'h2: w6aL01ok1NWMnhRdDAP = 32'd745594920 ^ 32'd2288768516 ^ 32'd2722199281;
      6'd7: w6aL01ok1NWMnhRdDAP = 32'b01010001111111011110100110100000 ^ 32'd1470605693;
      6'd31: w6aL01ok1NWMnhRdDAP = 32'd215854083 ^ 32'o7613363515 ^ 32'h34aa0b93;
      6'b110011: w6aL01ok1NWMnhRdDAP = 32'hf08014a8 ^ 32'd2175010107 ^ 32'b01110111011111100101000101001110;
      6'd17: w6aL01ok1NWMnhRdDAP = 32'd2827045785 ^ 32'd2933590852;
    endcase
  end

  logic [31:0] xQJVlE5Exe8992r1klC;
  always_comb begin
    case ({CLD6rGMxYQM8yZ4, raRSSx568gLgRd, C8sfwwEjm50H, LhC, jV8bIfqHdflwW, busy})
      6'd2: xQJVlE5Exe8992r1klC = 32'd3548693354 ^ 32'd3642768403;
      6'o1: xQJVlE5Exe8992r1klC = 32'b01111110000101010011001011111011 ^ 32'h211a156c ^ 32'h55abd8ef;
      6'b110011: xQJVlE5Exe8992r1klC = 32'b00100011000010001111011100011011 ^ 32'b00101001101011000000100001100010;
      6'd61: xQJVlE5Exe8992r1klC = 32'ha4780c4 ^ 32'b00000000111000110111111110111100;
      6'o73: xQJVlE5Exe8992r1klC = 32'd2679278382 ^ 32'o35725257042 ^ 32'o17220625165;
      6'o40: xQJVlE5Exe8992r1klC = 32'o22646243077 ^ 32'hb174e434 ^ 32'o5522256563;
      6'b110000: xQJVlE5Exe8992r1klC = 32'd284972748 ^ 32'h278a9e5f ^ 32'b00111101110100100011011111101011;
      6'o6: xQJVlE5Exe8992r1klC = 32'hccecb58d ^ 32'hc6484af4;
      6'h13: xQJVlE5Exe8992r1klC = 32'hc86d9773 ^ 32'b11011101001100110010110100101101 ^ 32'd536495399;
      6'b001100: xQJVlE5Exe8992r1klC = 32'h64eed518 ^ 32'b00000101111000000100011000010001 ^ 32'h6baa6c71;
      6'd16: xQJVlE5Exe8992r1klC = 32'd1584619500 ^ 32'd1423417492;
      6'b011111: xQJVlE5Exe8992r1klC = 32'b01011111110001100110000111100011 ^ 32'b01010101011000101001111010011010;
      6'o12: xQJVlE5Exe8992r1klC = 32'h6cfa0764 ^ 32'd1631002872 ^ 32'o732354345;
      6'b101000: xQJVlE5Exe8992r1klC = 32'd1968816295 ^ 32'b01111111111111010011111111011111;
      6'd38: xQJVlE5Exe8992r1klC = 32'b11011101011111111011010101001111 ^ 32'd1703789822 ^ 32'o26225507310;
      6'd35: xQJVlE5Exe8992r1klC = 32'ha6847e10 ^ 32'd1719455552 ^ 32'o31227047051;
      6'd55: xQJVlE5Exe8992r1klC = 32'd531442737 ^ 32'h1509d348;
      6'b010001: xQJVlE5Exe8992r1klC = 32'd1426243058 ^ 32'hc304d658 ^ 32'h9ca294d2;
      6'h39: xQJVlE5Exe8992r1klC = 32'o31260415631 ^ 32'h81d02d5e ^ 32'd1102498239;
      6'h0: xQJVlE5Exe8992r1klC = 32'b11011000011100000000100011011110 ^ 32'd124824826 ^ 32'b11010101101001000101101101011100;
      6'd22: xQJVlE5Exe8992r1klC = 32'he6369b26 ^ 32'd2011943430 ^ 32'b10011011011110011011011001011001;
      6'b001101: xQJVlE5Exe8992r1klC = 32'd690227189 ^ 32'b01011001110011110010000100011011 ^ 32'd2052053398;
      6'o3: xQJVlE5Exe8992r1klC = 32'h2d2744a5 ^ 32'o4740735734;
      6'd24: xQJVlE5Exe8992r1klC = 32'd1590834788 ^ 32'd1417070876;
      6'h8: xQJVlE5Exe8992r1klC = 32'hc242b251 ^ 32'd84127548 ^ 32'hcde5e215;
      6'b100100: xQJVlE5Exe8992r1klC = 32'o3531016511 ^ 32'd2490026464 ^ 32'b10000011101010100010101111010001;
      6'b010111: xQJVlE5Exe8992r1klC = 32'o24075514254 ^ 32'd2857527253;
      6'b000111: xQJVlE5Exe8992r1klC = 32'ha8f4bc21 ^ 32'o24224041530;
      6'd39: xQJVlE5Exe8992r1klC = 32'hc2277e61 ^ 32'd3364061464;
      6'b101011: xQJVlE5Exe8992r1klC = 32'he918fcea ^ 32'hb0cf41b1 ^ 32'o12334641042;
      6'd46: xQJVlE5Exe8992r1klC = 32'd3374300693 ^ 32'hc3bb416c;
      6'h1e: xQJVlE5Exe8992r1klC = 32'h501eb4e ^ 32'h746864a5 ^ 32'd2077061266;
      6'd27: xQJVlE5Exe8992r1klC = 32'o34575712404 ^ 32'd4015221373;
      6'o41: xQJVlE5Exe8992r1klC = 32'o12664656131 ^ 32'o13435721441;
      6'd52: xQJVlE5Exe8992r1klC = 32'd4096664028 ^ 32'd1511075173 ^ 32'd2761683905;
      6'd42: xQJVlE5Exe8992r1klC = 32'b10100010010010111111111001000000 ^ 32'o25073600471;
      6'b010100: xQJVlE5Exe8992r1klC = 32'b10101010000101110110110111110100 ^ 32'b01010111111111101100111111011010 ^ 32'o36723256526;
      6'b011101: xQJVlE5Exe8992r1klC = 32'hc51e0957 ^ 32'b11001111101110101111011000101111;
      6'd54: xQJVlE5Exe8992r1klC = 32'o35023471444 ^ 32'o34272506135;
      6'h29: xQJVlE5Exe8992r1klC = 32'd113385154 ^ 32'b00001100011001101110000110111010;
      6'o25: xQJVlE5Exe8992r1klC = 32'hf0a4f91c ^ 32'o37200003144;
      6'b100101: xQJVlE5Exe8992r1klC = 32'b10100010010010100010010101111000 ^ 32'h1a4d743f ^ 32'o26250727077;
      6'd60: xQJVlE5Exe8992r1klC = 32'h7aaaf999 ^ 32'hcb9ceb78 ^ 32'b10111011100100101110110110011001;
      6'o16: xQJVlE5Exe8992r1klC = 32'd2597524148 ^ 32'b00000101000000100001010001000100 ^ 32'h9575f989;
      6'b011010: xQJVlE5Exe8992r1klC = 32'd838867924 ^ 32'd950330541;
      6'd49: xQJVlE5Exe8992r1klC = 32'o6721524567 ^ 32'o7570453017;
      6'o77: xQJVlE5Exe8992r1klC = 32'd4123386271 ^ 32'b10111000011101010001101001110101 ^ 32'b01000111000101000000010010010011;
      6'b101111: xQJVlE5Exe8992r1klC = 32'heb98af41 ^ 32'd3571655725 ^ 32'o6567672025;
      6'b001111: xQJVlE5Exe8992r1klC = 32'h7cd48a66 ^ 32'o13511751313 ^ 32'o5325723724;
      6'd56: xQJVlE5Exe8992r1klC = 32'd2382335463 ^ 32'o20726671237;
      6'd11: xQJVlE5Exe8992r1klC = 32'd1229959180 ^ 32'h58471915 ^ 32'd464279136;
      6'h3e: xQJVlE5Exe8992r1klC = 32'o24336722302 ^ 32'o25167655673;
      6'b000101: xQJVlE5Exe8992r1klC = 32'o10066325123 ^ 32'd1249727787;
      6'h9: xQJVlE5Exe8992r1klC = 32'h4044a5b9 ^ 32'o11270055301;
      6'b101100: xQJVlE5Exe8992r1klC = 32'o20504503145 ^ 32'h7b47716e ^ 32'b11110100111100010000100001110011;
      6'h12: xQJVlE5Exe8992r1klC = 32'o27032143412 ^ 32'hb2cc3873;
      6'd28: xQJVlE5Exe8992r1klC = 32'b10101001110101011111001110010111 ^ 32'd2742095087;
      6'h32: xQJVlE5Exe8992r1klC = 32'h7cf344ba ^ 32'h7657bbc3;
      6'h2d: xQJVlE5Exe8992r1klC = 32'd2392889227 ^ 32'b11000000011001000000111100101100 ^ 32'h446067df;
      6'd34: xQJVlE5Exe8992r1klC = 32'd2775935452 ^ 32'b00110000011010010000011100111001 ^ 32'b10011111101110001001000110011100;
      6'd4: xQJVlE5Exe8992r1klC = 32'o27676651431 ^ 32'hb45fac61;
      6'o31: xQJVlE5Exe8992r1klC = 32'b00111101011111001011010110010001 ^ 32'o33344556476 ^ 32'o35422513727;
      6'h35: xQJVlE5Exe8992r1klC = 32'o36224071705 ^ 32'd2508668947 ^ 32'h6d73ccae;
      6'o72: xQJVlE5Exe8992r1klC = 32'b01001101001100100000001010010001 ^ 32'b01000111100101101111110111101000;
    endcase
  end

  always_ff @(posedge clk_i) begin
    if(rst_i) begin
      baudrate <= 9600;
    end else if (w6aL01ok1NWMnhRdDAP[32'h3cc51698 ^ 32'b00111100110001010001011010001000]) begin
      baudrate <= 9600;
    end else if(xQJVlE5Exe8992r1klC[32'o14647137617 ^ 32'h669cbf8f]) begin
      baudrate <= UIumLdEgx8;
    end
    else begin
      baudrate <= baudrate;
    end
  end

  logic WwX3PYk10uBYtDXg;
  assign WwX3PYk10uBYtDXg = UIumLdEgx8[32'b11000011111011111100010101000100 ^ 32'd3060869768 ^ 32'o16547567714];
  logic n3myOQv8Aqi;
  assign n3myOQv8Aqi = Pn7J == (32'd2842253610 ^ 32'ha969593a);
  logic [31:0] KleTBQQCTaG;

  always_comb begin
    case ({WwX3PYk10uBYtDXg, n3myOQv8Aqi, C8sfwwEjm50H, raRSSx568gLgRd, CLD6rGMxYQM8yZ4, LhC, parity_en})
      7'h3: KleTBQQCTaG = 32'h78d8d042 ^ 32'hbcb8004;
      7'b1110011: KleTBQQCTaG = 32'd2148291427 ^ 32'b11110011000111110000001100100101;
      7'd127: KleTBQQCTaG = 32'b10111010010000111011110000000000 ^ 32'h8950ec46;
      7'o51: KleTBQQCTaG = 32'o7207564613 ^ 32'h490db9cd;
      7'o145: KleTBQQCTaG = 32'h59488656 ^ 32'b00101010010110111101011000010000;
      7'h42: KleTBQQCTaG = 32'b01000110010010100111000010100101 ^ 32'ha8d822df ^ 32'o33540201074;
      7'ha: KleTBQQCTaG = 32'd2108675432 ^ 32'b01001110101111001000010100101110;
      7'd36: KleTBQQCTaG = 32'he226c268 ^ 32'o32115311056;
      7'h5e: KleTBQQCTaG = 32'd2803614861 ^ 32'd2018312738 ^ 32'b11101100010001011001011011101001;
      7'b1110101: KleTBQQCTaG = 32'h52d4330a ^ 32'd566715212;
      7'o120: KleTBQQCTaG = 32'd1400832814 ^ 32'h95db69f7 ^ 32'b11110101101101110011101010011111;
      7'o156: KleTBQQCTaG = 32'd3876964058 ^ 32'hd406969c;
      7'o144: KleTBQQCTaG = 32'b00111111011100111111011101001101 ^ 32'o15373607142 ^ 32'o14743724551;
      7'b0010010: KleTBQQCTaG = 32'h534fbaa7 ^ 32'b10010001100000001100011110111001 ^ 32'd4057738584;
      7'h5f: KleTBQQCTaG = 32'o3475354330 ^ 32'b10101000100001011111010111111111 ^ 32'd2271444321;
      7'd51: KleTBQQCTaG = 32'b10010010010100100100111010010011 ^ 32'd2715925263 ^ 32'b00000000101000001010010111011010;
      7'd76: KleTBQQCTaG = 32'b11111001100100000000100101010010 ^ 32'o6022224135 ^ 32'd4207571273;
      7'o142: KleTBQQCTaG = 32'b10100001111110010011011101111000 ^ 32'h92ea673e;
      7'o25: KleTBQQCTaG = 32'he7e22558 ^ 32'd4255233558 ^ 32'b01101001010100001100001100001000;
      7'o14: KleTBQQCTaG = 32'o16474422277 ^ 32'd2646301884 ^ 32'd3663341637;
      7'b1101100: KleTBQQCTaG = 32'hf9ed8e53 ^ 32'hcafede15;
      7'h60: KleTBQQCTaG = 32'o21051306567 ^ 32'b10111011101101101101110100110001;
      7'o126: KleTBQQCTaG = 32'h725511be ^ 32'd2185447366 ^ 32'd3271886398;
      7'd93: KleTBQQCTaG = 32'b00101111010001100100111100001101 ^ 32'hffe08466 ^ 32'ha3b59b2d;
      7'o74: KleTBQQCTaG = 32'h1c5006be ^ 32'b00101111010000110101011011111000;
      7'd59: KleTBQQCTaG = 32'o34233137305 ^ 32'o32137767203;
      7'd68: KleTBQQCTaG = 32'o31443350301 ^ 32'hc118ba85 ^ 32'b00111110100001100011101000000010;
      7'o10: KleTBQQCTaG = 32'b00110000000000011001110100110110 ^ 32'd51563888;
      7'h53: KleTBQQCTaG = 32'o14432045345 ^ 32'd393943715;
      7'b1011000: KleTBQQCTaG = 32'd1391492398 ^ 32'b01100001111000110010110101101000;
      7'b0100001: KleTBQQCTaG = 32'b11111100011110111111001110100101 ^ 32'h8f68a3e3;
      7'o107: KleTBQQCTaG = 32'o26154123734 ^ 32'o30250773632;
      7'h7b: KleTBQQCTaG = 32'd3751814289 ^ 32'b10101100101100110111010011010111;
      7'h7d: KleTBQQCTaG = 32'h4973fdab ^ 32'd1657676346 ^ 32'h58ae8fd7;
      7'o60: KleTBQQCTaG = 32'hd5de263e ^ 32'b11100110110011010111011001111000;
      7'd121: KleTBQQCTaG = 32'b00100011110100010010111101011100 ^ 32'h50c27f1a;
      7'h4b: KleTBQQCTaG = 32'b00011100001110111110000010000010 ^ 32'd3063599798 ^ 32'b11011001101100100110001001110010;
      7'o50: KleTBQQCTaG = 32'o33012160000 ^ 32'b11101011001110111011000001000110;
      7'd35: KleTBQQCTaG = 32'h341018b5 ^ 32'd3693510173 ^ 32'h9b2536ee;
      7'o76: KleTBQQCTaG = 32'b10011100100001101101110011011000 ^ 32'b10011100001100010011101000010101 ^ 32'd866432651;
      7'b0010011: KleTBQQCTaG = 32'd185230846 ^ 32'b01111000000110010011010110111000;
      7'h4a: KleTBQQCTaG = 32'o25001220655 ^ 32'b00101000011100000111110110011101 ^ 32'o26331406166;
      7'o13: KleTBQQCTaG = 32'h244f65fe ^ 32'b00100010001000010011010101000101 ^ 32'b01110101011111010000000011111101;
      7'o16: KleTBQQCTaG = 32'h99dedaf7 ^ 32'o34026562436 ^ 32'b01001010100101110110111110101111;
      7'h1: KleTBQQCTaG = 32'b11010110001001100101100110010011 ^ 32'b10001001011000001100001011011000 ^ 32'd743820045;
      7'o170: KleTBQQCTaG = 32'd1170600386 ^ 32'b01100101100110000000101011100001 ^ 32'd323922789;
      7'b1001101: KleTBQQCTaG = 32'o22003150754 ^ 32'b11100011000111111000000110101010;
      7'b0001111: KleTBQQCTaG = 32'o12373553461 ^ 32'b01100101101010110011000110001011 ^ 32'd1163310844;
      7'o53: KleTBQQCTaG = 32'h8af93c44 ^ 32'o37172466002;
      7'b0110010: KleTBQQCTaG = 32'd1634854689 ^ 32'd1382201191;
      7'o162: KleTBQQCTaG = 32'd4152116405 ^ 32'h846f14f3;
      7'o116: KleTBQQCTaG = 32'd1042194411 ^ 32'b00001101000011011100111110101101;
      7'd82: KleTBQQCTaG = 32'b00101000001010001100000001000101 ^ 32'd2055227391 ^ 32'd1639700476;
      7'o65: KleTBQQCTaG = 32'd1613448082 ^ 32'b10010011110100011010100101010000 ^ 32'b10000000111010011011101010000100;
      7'h45: KleTBQQCTaG = 32'b01100011011011110010000011010010 ^ 32'd276590740;
      7'h4: KleTBQQCTaG = 32'b10101110011010000101101111101000 ^ 32'o2715744241 ^ 32'o21223141417;
      7'd105: KleTBQQCTaG = 32'h3753a6b8 ^ 32'b00110101011101100100110110010001 ^ 32'd1899412335;
      7'h1b: KleTBQQCTaG = 32'd2270272602 ^ 32'b00101100011110101110110110010001 ^ 32'o33016020615;
      7'b1101011: KleTBQQCTaG = 32'o25757106451 ^ 32'b01111101001001110000111110101010 ^ 32'o24142151305;
      7'd111: KleTBQQCTaG = 32'b01101001001001111000110000000100 ^ 32'b00011010001101001101110001000010;
      7'b0000010: KleTBQQCTaG = 32'o24044767000 ^ 32'o12066606262 ^ 32'o30326731364;
      7'o132: KleTBQQCTaG = 32'o21056776771 ^ 32'o31156022651 ^ 32'b01110010000100001000100000010110;
      7'h34: KleTBQQCTaG = 32'b00100100010101010111010011101100 ^ 32'd3543223875 ^ 32'd3296160489;
      7'h14: KleTBQQCTaG = 32'd2561999675 ^ 32'o25351451575;
      7'b1010111: KleTBQQCTaG = 32'b01100000100001010001011010111101 ^ 32'ha2e9a361 ^ 32'o26137762632;
      7'b1100001: KleTBQQCTaG = 32'd2337084233 ^ 32'h7bb50be1 ^ 32'd2213234926;
      7'd102: KleTBQQCTaG = 32'h6f77ab36 ^ 32'b10010011101110111001011101101101 ^ 32'hcfdf6c1d;
      7'o46: KleTBQQCTaG = 32'd2822831856 ^ 32'habafa8a6 ^ 32'b00110000111111000000011000010000;
      7'd89: KleTBQQCTaG = 32'hbcbcb456 ^ 32'h4df65e38 ^ 32'h8259ba28;
      7'o52: KleTBQQCTaG = 32'h8a6d893b ^ 32'h1d377f3b ^ 32'd2756290118;
      7'h6d: KleTBQQCTaG = 32'o14701636662 ^ 32'b00101000100101001110011111111101 ^ 32'o7440105011;
      7'o54: KleTBQQCTaG = 32'b10100010000011001010010011011011 ^ 32'd2434790557;
      7'd119: KleTBQQCTaG = 32'hf0fa1be0 ^ 32'd2213104550;
      7'o56: KleTBQQCTaG = 32'hb64aa2b7 ^ 32'b10000101010110011111001011110001;
      7'h1c: KleTBQQCTaG = 32'o22614263235 ^ 32'h7c26bf13 ^ 32'd3640953288;
      7'd124: KleTBQQCTaG = 32'b11101110100000100000001100011110 ^ 32'b10000101111101011110111000111000 ^ 32'o13031136540;
      7'd65: KleTBQQCTaG = 32'b01001101000100111110000100110111 ^ 32'b00111110000000001011000101110001;
      7'b0000000: KleTBQQCTaG = 32'b10111110111111110111010110010101 ^ 32'o23645357235 ^ 32'd326761294;
      7'o111: KleTBQQCTaG = 32'ha11ae053 ^ 32'b00111010000001001000001011111101 ^ 32'd3893179112;
      7'o26: KleTBQQCTaG = 32'b01000110111011110110110000001100 ^ 32'b01110101111111000011110001001010;
      7'd56: KleTBQQCTaG = 32'b00110100110000110010100000011101 ^ 32'h7d0785b;
      7'b1101000: KleTBQQCTaG = 32'o4554777336 ^ 32'd379629208;
      7'd29: KleTBQQCTaG = 32'hfbe3cd25 ^ 32'b11110010101101011110110100010100 ^ 32'd2051371127;
      7'o152: KleTBQQCTaG = 32'o6132656406 ^ 32'b00000010011110000000110101000000;
      7'd39: KleTBQQCTaG = 32'o12113762137 ^ 32'd574403609;
      7'o36: KleTBQQCTaG = 32'd3132637026 ^ 32'd2309713700;
      7'h3d: KleTBQQCTaG = 32'hb421f932 ^ 32'o30714524564;
      7'd70: KleTBQQCTaG = 32'd3759102312 ^ 32'b11010011000111000000100100101110;
      7'b0010000: KleTBQQCTaG = 32'b00000111000110000000101001001000 ^ 32'b11001010111000001011010001110010 ^ 32'o37672767174;
      7'hd: KleTBQQCTaG = 32'o34055663416 ^ 32'd1238909636 ^ 32'b11011010011111000111010110001100;
      7'd26: KleTBQQCTaG = 32'o15541107202 ^ 32'o13645757304;
      7'd31: KleTBQQCTaG = 32'b01001001010010110101001110010011 ^ 32'o11210464034 ^ 32'd813329353;
      7'd99: KleTBQQCTaG = 32'b11111000001111101010111101010000 ^ 32'o2113171145 ^ 32'd2583760243;
      7'b0010111: KleTBQQCTaG = 32'b10101110100101001111000100110001 ^ 32'b11011101100001111010000101110111;
      7'd122: KleTBQQCTaG = 32'b00101010111100010100101001001111 ^ 32'd809425953 ^ 32'o15167143050;
      7'd112: KleTBQQCTaG = 32'o24351310706 ^ 32'o22055540600;
      7'b1011100: KleTBQQCTaG = 32'd1434699467 ^ 32'b01100110100100001001011010001101;
      7'd57: KleTBQQCTaG = 32'd3832947299 ^ 32'd2241702071 ^ 32'b00010010111110001101101010010010;
      7'd84: KleTBQQCTaG = 32'h65b161c5 ^ 32'o33705417453 ^ 32'd2310287016;
      7'd17: KleTBQQCTaG = 32'd204905259 ^ 32'd2133183341;
      7'd7: KleTBQQCTaG = 32'd1392021155 ^ 32'd3587981614 ^ 32'b11110100001101111001111111001011;
      7'd9: KleTBQQCTaG = 32'd3433211555 ^ 32'hbfb1f6e5;
      7'b0011001: KleTBQQCTaG = 32'h2f666397 ^ 32'd2487279357 ^ 32'o31015366454;
      7'b1000000: KleTBQQCTaG = 32'd119959048 ^ 32'd875904590;
      7'b0101111: KleTBQQCTaG = 32'hc40d625 ^ 32'd2136180323;
      7'b0110110: KleTBQQCTaG = 32'b11001111001010000101111000111001 ^ 32'b11111100001110110000111001111111;
      7'b0110001: KleTBQQCTaG = 32'b00001101110000100011001001000010 ^ 32'h7ed16204;
      7'b1111110: KleTBQQCTaG = 32'd2973985533 ^ 32'h82503abb;
      7'b1011011: KleTBQQCTaG = 32'o17662400306 ^ 32'o1566250200;
      7'h22: KleTBQQCTaG = 32'd1873282540 ^ 32'b01001101111111000001010110101010 ^ 32'b00010001010001110100000000000000;
      7'o110: KleTBQQCTaG = 32'd4272280305 ^ 32'd3451290295;
      7'o45: KleTBQQCTaG = 32'd1060508817 ^ 32'h8aac0c84 ^ 32'o30642244123;
      7'b1100111: KleTBQQCTaG = 32'b01010010110010011110111011111111 ^ 32'b00100001110110101011111010111001;
      7'd81: KleTBQQCTaG = 32'o13627302612 ^ 32'h2d4ed5cc;
      7'd24: KleTBQQCTaG = 32'hf005a13c ^ 32'b11000011000101101111000101111010;
      7'b1110001: KleTBQQCTaG = 32'o35342435320 ^ 32'd2560191126;
      7'd58: KleTBQQCTaG = 32'b01011010110010111110111000000001 ^ 32'o27266711335 ^ 32'b11010011000000110010110010011010;
      7'b1110110: KleTBQQCTaG = 32'd1416661077 ^ 32'o4730754023;
      7'h55: KleTBQQCTaG = 32'd1505420482 ^ 32'd715764868;
      7'o55: KleTBQQCTaG = 32'o32361347162 ^ 32'ha0d69e34;
      7'o103: KleTBQQCTaG = 32'd2754053393 ^ 32'd3212196731 ^ 32'd1749216812;
      7'h6: KleTBQQCTaG = 32'h99dfab26 ^ 32'b10101010110011001111101101100000;
      7'o77: KleTBQQCTaG = 32'o30273675245 ^ 32'b11110001111111000010101011100011;
      7'o40: KleTBQQCTaG = 32'hed8e3e1c ^ 32'o33647267132;
      7'b0000101: KleTBQQCTaG = 32'o21342544110 ^ 32'b11000110110001100101000010111011 ^ 32'd1046464693;
      7'd55: KleTBQQCTaG = 32'haa3dc4d2 ^ 32'h1532440a ^ 32'b10001100000111001101000010011110;
      7'o117: KleTBQQCTaG = 32'h7191ee39 ^ 32'h282be7f;
      7'o164: KleTBQQCTaG = 32'o34311725332 ^ 32'h6bf5ba95 ^ 32'b10111011110000010100000000001001;
    endcase
  end

  always_ff @(posedge clk_i) begin
    if(rst_i) begin
      parity_en <= '0;
    end
    else begin
      parity_en <= KleTBQQCTaG[32'o15162645033 ^ 32'd2306009849 ^ 32'he0b9a0fc];
    end
  end

  logic i16aOBIRoTka;
  assign i16aOBIRoTka = Pn7J == (32'h5dd503ee ^ 32'o33420446676 ^ 32'd2174176836);

  logic [31:0] cwp;
  logic [31:0] aboba;

  always_comb begin
    case ({i16aOBIRoTka, raRSSx568gLgRd, C8sfwwEjm50H, CLD6rGMxYQM8yZ4, LhC})
      5'd20: cwp = 32'b00010010111100100100110111100001 ^ 32'hfb0489a;
      5'o4: cwp = 32'hf4f8aa0b ^ 32'd3921325936;
      5'b00001: cwp = 32'o13052166122 ^ 32'h45eae929;
      5'h16: cwp = 32'ha35e7b3f ^ 32'hbe1c7e44;
      5'd5: cwp = 32'd2888127131 ^ 32'h40fd1d16 ^ 32'd4053420790;
      5'b11111: cwp = 32'h7a45cc3 ^ 32'o12215157665 ^ 32'h48c2860d;
      5'b11010: cwp = 32'o34234343312 ^ 32'o37714741661;
      5'd13: cwp = 32'd4221104830 ^ 32'd2340652064 ^ 32'o15526271745;
      5'd28: cwp = 32'd2432621365 ^ 32'hae340fd ^ 32'd2271190707;
      5'he: cwp = 32'o12545735456 ^ 32'b10111011101000010010101110010011 ^ 32'b11110011011101001001010111000110;
      5'h11: cwp = 32'o7553445060 ^ 32'o4073047513;
      5'd8: cwp = 32'b11010010011000001001101111001110 ^ 32'o31710517265;
      5'd16: cwp = 32'b10000111010100111110000001110000 ^ 32'o21774000510 ^ 32'o2570362103;
      5'b11110: cwp = 32'ha60cd27d ^ 32'd3142506246;
      5'ha: cwp = 32'b11011011101001000001101100001011 ^ 32'o30671417160;
      5'd29: cwp = 32'd2027720029 ^ 32'b01101010101000000111100010111000 ^ 32'hf3ef09e;
      5'o17: cwp = 32'h478b12da ^ 32'b00111111000111000011110000011100 ^ 32'o14561225675;
      5'h6: cwp = 32'b10011110011100101100001010010001 ^ 32'b10000011001100001100011111101010;
      5'h7: cwp = 32'd1052590111 ^ 32'h23ff4564;
      5'b11011: cwp = 32'b11110000010100100101010010100000 ^ 32'h6262e94 ^ 32'd3946217295;
      5'd3: cwp = 32'b01000110011000001010000001011111 ^ 32'b01011011001000101010010100100100;
      5'd11: cwp = 32'ha8d7ede1 ^ 32'd3046500506;
      5'd12: cwp = 32'b01111000100101010000011011000101 ^ 32'b11001101100001101000111110011010 ^ 32'o25024306044;
      5'h15: cwp = 32'd2664618246 ^ 32'b10000011100100001101110001111101;
      5'o27: cwp = 32'd3691529365 ^ 32'd3242869230;
      5'o0: cwp = 32'o5427444531 ^ 32'd823938082;
      5'b01001: cwp = 32'o2371101674 ^ 32'd1222139078 ^ 32'o10637555001;
      5'd24: cwp = 32'h4f54efea ^ 32'o35157175344 ^ 32'd3148484725;
      5'o2: cwp = 32'o32343615617 ^ 32'b11001110110011010001111011110100;
      5'd19: cwp = 32'b01100101010000000000110011011011 ^ 32'b01111000000000100000100110100000;
      5'h12: cwp = 32'b10000000100011111001111011111001 ^ 32'h52f26fee ^ 32'o31717772154;
      5'd25: cwp = 32'had7dde7a ^ 32'o26017755401;
      default: cwp = 32'hdead_dead;
    endcase
  end

  assign       l4fxxX4aa = Pn7J == (32'hce2043db ^ 32'b00010101000100111011110101010100 ^ 32'b11011011001100111111111010000111);

  always_ff @(posedge clk_i) begin
    if(rst_i) begin
      stopbit <= '0;
    end
    else if (cwp[32'd1173052495 ^ 32'h45eb5c5b]) begin
      stopbit <= '0;
    end
    else if(aboba[32'b10001101000100111101110110111101 ^ 32'b10001101000100111101110110111101]) begin
      stopbit <= UIumLdEgx8[1:0];
    end
    else begin
      stopbit <= stopbit;
    end
  end
  assign jV8bIfqHdflwW = Pn7J == (32'd1055356197 ^ 32'd1055356201);

  always_comb begin
    case ({i16aOBIRoTka, raRSSx568gLgRd, C8sfwwEjm50H, CLD6rGMxYQM8yZ4, LhC})
      5'ha: aboba = 32'h3087f3dc ^ 32'o10402636570;
      5'b00101: aboba = 32'h271e5554 ^ 32'b11111001011001100110101001001000 ^ 32'haaf4f1b8;
      5'o34: aboba = 32'd849669163 ^ 32'o10334524566 ^ 32'o526505771;
      5'b01111: aboba = 32'b11110101011110010100000001100101 ^ 32'd3044917641 ^ 32'b00110100100010000100111101001000;
      5'o22: aboba = 32'b11010101001111101000011000010011 ^ 32'h87bb5ecd ^ 32'd638129786;
      5'o23: aboba = 32'b11001000001011000000100001011101 ^ 32'd4094572533 ^ 32'd1219424524;
      5'o32: aboba = 32'd811175085 ^ 32'b10100010001010111100000111100000 ^ 32'he6fe83e9;
      5'b00011: aboba = 32'o34053244436 ^ 32'd595348521 ^ 32'hb75dcb93;
      5'b00110: aboba = 32'd3776296783 ^ 32'b01110101010000010000000001101100 ^ 32'd3772283271;
      5'b00100: aboba = 32'd810798815 ^ 32'd1155465339;
      5'o25: aboba = 32'd1585867373 ^ 32'o5202522310;
      5'o20: aboba = 32'he3230c2b ^ 32'd3308654975 ^ 32'b01010010100110011101001111110000;
      5'b00000: aboba = 32'o34677371106 ^ 32'b01110111010110001110000001010110 ^ 32'd3844725940;
      5'b01101: aboba = 32'h53fbbbb3 ^ 32'd662140183;
      5'b11000: aboba = 32'b10000001100111111110110010001110 ^ 32'o1744525771 ^ 32'hfa8189d3;
      5'he: aboba = 32'd2876869146 ^ 32'd3892100178 ^ 32'o7002374354;
      5'h19: aboba = 32'd3671789667 ^ 32'h7d2ec349 ^ 32'hd3791d8e;
      5'o21: aboba = 32'h1201096a ^ 32'b01100110100011011100011111001110;
      5'h9: aboba = 32'hf1d03daa ^ 32'd2237461262;
      5'o14: aboba = 32'd306409911 ^ 32'o14663737423;
      5'b10110: aboba = 32'b01000000011111110110010010011010 ^ 32'd888384062;
      5'b11101: aboba = 32'b01111000000110111010010011000101 ^ 32'o1445665140;
      5'h7: aboba = 32'hd87c8880 ^ 32'o11776070274 ^ 32'o34302033230;
      5'h1b: aboba = 32'hbbede754 ^ 32'o24534230725 ^ 32'o15204014045;
      5'h1e: aboba = 32'd4063396739 ^ 32'o20657446447;
      5'd20: aboba = 32'd682760427 ^ 32'h5c3ed64f;
      5'o10: aboba = 32'd1917169571 ^ 32'd113860871;
      5'hb: aboba = 32'b01101110100011001011001010000000 ^ 32'h1a007c24;
      5'h2: aboba = 32'd2792801143 ^ 32'd3539602899;
      5'h1: aboba = 32'd2135621536 ^ 32'b10001101010010110110011101101111 ^ 32'o20643253153;
      5'b11111: aboba = 32'o24323057554 ^ 32'h3825728e ^ 32'd4024820551;
      5'b10111: aboba = 32'd2427150063 ^ 32'o34042706360 ^ 32'o453016272;
      default: aboba = 32'hdead_dead;
    endcase
  end

  always_comb begin
    case ({raRSSx568gLgRd, C8sfwwEjm50H, LhC, WwX3PYk10uBYtDXg, CLD6rGMxYQM8yZ4})
      5'h1c: cSJpl8RGMw2bgs48nEfg = 32'd2048862294 ^ 32'b10111001011101111101011011001001 ^ 32'h89ab6b30;
      5'o1: cSJpl8RGMw2bgs48nEfg = 32'h4702ec71 ^ 32'h9e3dcd92 ^ 32'b10010011111111001011010001001100;
      5'hf: cSJpl8RGMw2bgs48nEfg = 32'b10011111000000011010010001001000 ^ 32'o32560430747;
      5'b11000: cSJpl8RGMw2bgs48nEfg = 32'b10001010111010011100010110101111 ^ 32'd142793182 ^ 32'o31052104736;
      5'h15: cSJpl8RGMw2bgs48nEfg = 32'd2470939058 ^ 32'o21043235574 ^ 32'b01010001000010010010011101100001;
      5'd6: cSJpl8RGMw2bgs48nEfg = 32'b11000100111110110100011101010100 ^ 32'd2386088699;
      5'o20: cSJpl8RGMw2bgs48nEfg = 32'b10100000111101010100110011111110 ^ 32'b11101010001101101101100101010001;
      5'd11: cSJpl8RGMw2bgs48nEfg = 32'hcea947bb ^ 32'b10100110000111110100001010001001 ^ 32'h2275909d;
      5'b11111: cSJpl8RGMw2bgs48nEfg = 32'b01100000011001001001011010001100 ^ 32'd715326243;
      5'd10: cSJpl8RGMw2bgs48nEfg = 32'd2041134147 ^ 32'h336aa9ec;
      5'h19: cSJpl8RGMw2bgs48nEfg = 32'o1014251566 ^ 32'o21534247460 ^ 32'd3481504233;
      5'd2: cSJpl8RGMw2bgs48nEfg = 32'hfc763156 ^ 32'hb6b5a4f9;
      5'b00111: cSJpl8RGMw2bgs48nEfg = 32'b01000010010010000011001011111111 ^ 32'b11100111110111000101011010011111 ^ 32'd4015518159;
      5'o15: cSJpl8RGMw2bgs48nEfg = 32'b01001110000011011001111110000110 ^ 32'h4ce0a29;
      5'd17: cSJpl8RGMw2bgs48nEfg = 32'd3953211026 ^ 32'h644ea49c ^ 32'b11000101001011000000011110100001;
      5'b01000: cSJpl8RGMw2bgs48nEfg = 32'd779271157 ^ 32'b01100100101100010010111001011010;
      5'd12: cSJpl8RGMw2bgs48nEfg = 32'o36075552706 ^ 32'hd4aa6d79 ^ 32'b01101110100111110010110100010000;
      5'd4: cSJpl8RGMw2bgs48nEfg = 32'b11011111101101000100110101110010 ^ 32'o22535754335;
      5'o24: cSJpl8RGMw2bgs48nEfg = 32'd1010024144 ^ 32'hbb72f903 ^ 32'b11001101100000101101001001111100;
      5'b10011: cSJpl8RGMw2bgs48nEfg = 32'h2823d952 ^ 32'hb9b94f1a ^ 32'd3680044007;
      5'o5: cSJpl8RGMw2bgs48nEfg = 32'b10110011001110001001001000011101 ^ 32'b11111001111110110000011110110010;
      5'o27: cSJpl8RGMw2bgs48nEfg = 32'd2464334183 ^ 32'haf3a04db ^ 32'o16706650023;
      5'o33: cSJpl8RGMw2bgs48nEfg = 32'hd0593c12 ^ 32'h9a9aa9bd;
      5'h1d: cSJpl8RGMw2bgs48nEfg = 32'b10011001010101010111000111000110 ^ 32'd140435213 ^ 32'hdbcc3b64;
      5'd26: cSJpl8RGMw2bgs48nEfg = 32'h1daefd78 ^ 32'd1466788055;
      5'd9: cSJpl8RGMw2bgs48nEfg = 32'o565171552 ^ 32'h4f1766c5;
      5'o16: cSJpl8RGMw2bgs48nEfg = 32'hf3444dc5 ^ 32'd3681802092 ^ 32'd1660161798;
      5'd22: cSJpl8RGMw2bgs48nEfg = 32'he68f96ee ^ 32'b11011100010011101000011001101100 ^ 32'o16000502455;
      5'b00000: cSJpl8RGMw2bgs48nEfg = 32'hff840b1c ^ 32'o34604310746 ^ 32'd1398148949;
      5'b11110: cSJpl8RGMw2bgs48nEfg = 32'hf3336a00 ^ 32'b10111001111100001111111110101111;
      5'h12: cSJpl8RGMw2bgs48nEfg = 32'o10321063242 ^ 32'b01000011011101000111000000010011 ^ 32'o11274701436;
      5'h3: cSJpl8RGMw2bgs48nEfg = 32'o36756405077 ^ 32'b10111101011110011001111110010000;
    endcase
  end

  always_comb begin
    case ({CLD6rGMxYQM8yZ4, LhC, WwX3PYk10uBYtDXg, C8sfwwEjm50H, raRSSx568gLgRd})
      5'd2: dNVOskLQGaCf26HqGY = 32'b11001111101011101101110001010111 ^ 32'h843e6b86;
      5'h19: dNVOskLQGaCf26HqGY = 32'hf9a82f7f ^ 32'o26216114252;
      5'h10: dNVOskLQGaCf26HqGY = 32'o10333464617 ^ 32'h8fede5e;
      5'b10111: dNVOskLQGaCf26HqGY = 32'd1352730113 ^ 32'o3314330720;
      5'd12: dNVOskLQGaCf26HqGY = 32'o34044007753 ^ 32'b01100011011100100110101100011001 ^ 32'b11001000011100101101001100100111;
      5'd5: dNVOskLQGaCf26HqGY = 32'o26642015215 ^ 32'o37506126534;
      5'b11100: dNVOskLQGaCf26HqGY = 32'h596a8671 ^ 32'd421143133 ^ 32'd199234553;
      5'h1: dNVOskLQGaCf26HqGY = 32'b11001111111101001010000010111010 ^ 32'b01110110001111111111001000001011 ^ 32'hf25be560;
      5'd4: dNVOskLQGaCf26HqGY = 32'b10010000100100111010000001000111 ^ 32'd3674412950;
      5'h1d: dNVOskLQGaCf26HqGY = 32'd1768120639 ^ 32'b00100010111100111101011011101010;
      5'o0: dNVOskLQGaCf26HqGY = 32'o23715253332 ^ 32'd3836222473 ^ 32'b00110000000011011111110100000010;
      5'h9: dNVOskLQGaCf26HqGY = 32'b00011101001101111000010001110101 ^ 32'h56a733a0;
      5'o3: dNVOskLQGaCf26HqGY = 32'o24576132517 ^ 32'd3999793822;
      5'd7: dNVOskLQGaCf26HqGY = 32'd3160163318 ^ 32'h58751096 ^ 32'o25756362261;
      5'o12: dNVOskLQGaCf26HqGY = 32'h6818fdce ^ 32'h8b72601e ^ 32'ha8fa2a01;
      5'b10101: dNVOskLQGaCf26HqGY = 32'hb2c420e7 ^ 32'hf9549736;
      5'o22: dNVOskLQGaCf26HqGY = 32'o12374714233 ^ 32'b00011000011000110010111101001010;
      5'b11111: dNVOskLQGaCf26HqGY = 32'hc38c6640 ^ 32'h881cd191;
      5'h1e: dNVOskLQGaCf26HqGY = 32'd1405343188 ^ 32'd408117765;
      5'o26: dNVOskLQGaCf26HqGY = 32'o35321477447 ^ 32'b11100111111000001011111110110100 ^ 32'h47367742;
      5'hf: dNVOskLQGaCf26HqGY = 32'b01011111000110000001010011110110 ^ 32'h1488a327;
      5'h6: dNVOskLQGaCf26HqGY = 32'o20676724556 ^ 32'd3446349503;
      5'h13: dNVOskLQGaCf26HqGY = 32'hd14592d8 ^ 32'd2125539496 ^ 32'he4640da1;
      5'o15: dNVOskLQGaCf26HqGY = 32'b00100010010101001110010110010001 ^ 32'o15161051104;
      5'b10100: dNVOskLQGaCf26HqGY = 32'o14572510074 ^ 32'b00101110110111111110100111101101 ^ 32'o51347000;
      5'o13: dNVOskLQGaCf26HqGY = 32'h7d7bb931 ^ 32'o6672607340;
      5'o10: dNVOskLQGaCf26HqGY = 32'b00010110101001001101111100101110 ^ 32'h708636c6 ^ 32'o5554457075;
      5'b10001: dNVOskLQGaCf26HqGY = 32'o32032450626 ^ 32'd3222387735 ^ 32'b01011011111010110101101001010000;
      5'h18: dNVOskLQGaCf26HqGY = 32'hee37065e ^ 32'b10100101101001111011000110001011;
      5'd27: dNVOskLQGaCf26HqGY = 32'h477b8ae6 ^ 32'h734d4e09 ^ 32'o17751471476;
      5'o32: dNVOskLQGaCf26HqGY = 32'd539038598 ^ 32'd64536488 ^ 32'd1751718911;
      5'he: dNVOskLQGaCf26HqGY = 32'h26f1bd77 ^ 32'ha48f1219 ^ 32'hc9ee18bf;
    endcase
  end
endmodule
