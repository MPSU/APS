module led_sb_ctrl(
/*
    Часть интерфейса модуля, отвечающая за подключение к системной шине
*/
  input  logic        clk_i,
  input  logic        rst_i,
  input  logic        req_i,
  input  logic        write_enable_i,
  input  logic [31:0] addr_i,
  input  logic [31:0] write_data_i,
  output logic [31:0] read_data_o,

/*
    Часть интерфейса модуля, отвечающая за подключение к периферии
*/
  output logic [15:0]  led_o
);
logic [15:0]  led_val;
logic         led_mode;

logic [31:0]  cntr;

logic soft_reset;

logic  soft_reset_addr_cmp;
assign soft_reset_addr_cmp = addr_i == 32'h24;

logic  soft_reset_write_data_cmp;
assign soft_reset_write_data_cmp = write_data_i == 1'b1;

assign soft_reset = req_i & write_enable_i & soft_reset_addr_cmp & soft_reset_write_data_cmp;

assign led_o = cntr < 32'd10_000_000 ? led_val : 32'd0;

logic  led_mode_addr_cmp;
assign led_mode_addr_cmp = addr_i == 32'd4;

logic  led_mode_write_data_cmp;
assign led_mode_write_data_cmp = write_data_i <= 32'd1;

logic led_mode_en;
always_comb begin
  case ({soft_reset_addr_cmp, led_mode_write_data_cmp, led_mode_addr_cmp, write_enable_i, req_i, soft_reset_write_data_cmp})
    6'b000000: led_mode_en = 1'b0;
    6'b000001: led_mode_en = 1'b0;
    6'b000010: led_mode_en = 1'b0;
    6'b000011: led_mode_en = 1'b0;
    6'b000100: led_mode_en = 1'b0;
    6'b000101: led_mode_en = 1'b0;
    6'b000110: led_mode_en = 1'b0;
    6'b000111: led_mode_en = 1'b0;
    6'b001000: led_mode_en = 1'b0;
    6'b001001: led_mode_en = 1'b0;
    6'b001010: led_mode_en = 1'b0;
    6'b001011: led_mode_en = 1'b0;
    6'b001100: led_mode_en = 1'b0;
    6'b001101: led_mode_en = 1'b0;
    6'b001110: led_mode_en = 1'b0;
    6'b001111: led_mode_en = 1'b0;
    6'b010000: led_mode_en = 1'b0;
    6'b010001: led_mode_en = 1'b0;
    6'b010010: led_mode_en = 1'b0;
    6'b010011: led_mode_en = 1'b0;
    6'b010100: led_mode_en = 1'b0;
    6'b010101: led_mode_en = 1'b0;
    6'b010110: led_mode_en = 1'b0;
    6'b010111: led_mode_en = 1'b0;
    6'b011000: led_mode_en = 1'b0;
    6'b011001: led_mode_en = 1'b0;
    6'b011010: led_mode_en = 1'b0;
    6'b011011: led_mode_en = 1'b0;
    6'b011100: led_mode_en = 1'b0;
    6'b011101: led_mode_en = 1'b0;
    6'b011110: led_mode_en = 1'b1;
    6'b011111: led_mode_en = 1'b1;
    6'b100000: led_mode_en = 1'b0;
    6'b100001: led_mode_en = 1'b0;
    6'b100010: led_mode_en = 1'b0;
    6'b100011: led_mode_en = 1'b0;
    6'b100100: led_mode_en = 1'b0;
    6'b100101: led_mode_en = 1'b0;
    6'b100110: led_mode_en = 1'b0;
    6'b100111: led_mode_en = 1'b1; // reset
    6'b101000: led_mode_en = 1'b0;
    6'b101001: led_mode_en = 1'b0;
    6'b101010: led_mode_en = 1'b0;
    6'b101011: led_mode_en = 1'b0;
    6'b101100: led_mode_en = 1'b0;
    6'b101101: led_mode_en = 1'b0;
    6'b101110: led_mode_en = 1'b0;
    6'b101111: led_mode_en = 1'b1; // reset
    6'b110000: led_mode_en = 1'b0;
    6'b110001: led_mode_en = 1'b0;
    6'b110010: led_mode_en = 1'b0;
    6'b110011: led_mode_en = 1'b0;
    6'b110100: led_mode_en = 1'b0;
    6'b110101: led_mode_en = 1'b0;
    6'b110110: led_mode_en = 1'b0;
    6'b110111: led_mode_en = 1'b1; // reset
    6'b111000: led_mode_en = 1'b0;
    6'b111001: led_mode_en = 1'b0;
    6'b111010: led_mode_en = 1'b0;
    6'b111011: led_mode_en = 1'b0;
    6'b111100: led_mode_en = 1'b0;
    6'b111101: led_mode_en = 1'b0;
    6'b111110: led_mode_en = 1'b1;
    6'b111111: led_mode_en = 1'b1; // reset
  endcase
end

logic  led_mode_next;
always_comb begin
  case ({req_i, write_data_i[0], write_enable_i, soft_reset_addr_cmp, soft_reset_write_data_cmp})
    5'b00000: led_mode_next = 1'b0;
    5'b00001: led_mode_next = 1'b0;
    5'b00010: led_mode_next = 1'b0;
    5'b00011: led_mode_next = 1'b0;
    5'b00100: led_mode_next = 1'b0;
    5'b00101: led_mode_next = 1'b0;
    5'b00110: led_mode_next = 1'b0;
    5'b00111: led_mode_next = 1'b0;
    5'b01000: led_mode_next = 1'b1;
    5'b01001: led_mode_next = 1'b1;
    5'b01010: led_mode_next = 1'b1;
    5'b01011: led_mode_next = 1'b1;
    5'b01100: led_mode_next = 1'b1;
    5'b01101: led_mode_next = 1'b1;
    5'b01110: led_mode_next = 1'b1;
    5'b01111: led_mode_next = 1'b1;
    5'b10000: led_mode_next = 1'b0;
    5'b10001: led_mode_next = 1'b0;
    5'b10010: led_mode_next = 1'b0;
    5'b10011: led_mode_next = 1'b0;
    5'b10100: led_mode_next = 1'b0;
    5'b10101: led_mode_next = 1'b0;
    5'b10110: led_mode_next = 1'b0;
    5'b10111: led_mode_next = 1'b0; // reset
    5'b11000: led_mode_next = 1'b1;
    5'b11001: led_mode_next = 1'b1;
    5'b11010: led_mode_next = 1'b1;
    5'b11011: led_mode_next = 1'b1;
    5'b11100: led_mode_next = 1'b1;
    5'b11101: led_mode_next = 1'b1;
    5'b11110: led_mode_next = 1'b1;
    5'b11111: led_mode_next = 1'b0; // reset
  endcase
end

always_ff @(posedge clk_i) begin
  if(rst_i) begin
    led_mode <= 1'b0;
  end else if(led_mode_en) begin
    led_mode <= led_mode_next;
  end
end

logic  cntr_cmp;
assign cntr_cmp = cntr < 32'd20_000_000;

logic [31:0] cntr_next;
always_comb begin
  case ({cntr_cmp, req_i, write_enable_i, soft_reset_addr_cmp, led_mode, soft_reset_write_data_cmp})
    6'b000000: cntr_next = '0;
    6'b000001: cntr_next = '0;
    6'b000010: cntr_next = '0;
    6'b000011: cntr_next = '0;
    6'b000100: cntr_next = '0;
    6'b000101: cntr_next = '0;
    6'b000110: cntr_next = '0;
    6'b000111: cntr_next = '0;
    6'b001000: cntr_next = '0;
    6'b001001: cntr_next = '0;
    6'b001010: cntr_next = '0;
    6'b001011: cntr_next = '0;
    6'b001100: cntr_next = '0;
    6'b001101: cntr_next = '0;
    6'b001110: cntr_next = '0;
    6'b001111: cntr_next = '0;
    6'b010000: cntr_next = '0;
    6'b010001: cntr_next = '0;
    6'b010010: cntr_next = '0;
    6'b010011: cntr_next = '0;
    6'b010100: cntr_next = '0;
    6'b010101: cntr_next = '0;
    6'b010110: cntr_next = '0;
    6'b010111: cntr_next = '0;
    6'b011000: cntr_next = '0;
    6'b011001: cntr_next = '0;
    6'b011010: cntr_next = '0;
    6'b011011: cntr_next = '0;
    6'b011100: cntr_next = '0;
    6'b011101: cntr_next = '0; // reset
    6'b011110: cntr_next = '0;
    6'b011111: cntr_next = '0; // reset

    6'b100000: cntr_next = '0;
    6'b100001: cntr_next = '0;
    6'b100010: cntr_next = cntr + 32'b1;
    6'b100011: cntr_next = cntr + 32'b1;
    6'b100100: cntr_next = '0;
    6'b100101: cntr_next = '0;
    6'b100110: cntr_next = cntr + 32'b1;
    6'b100111: cntr_next = cntr + 32'b1;
    6'b101000: cntr_next = '0;
    6'b101001: cntr_next = '0;
    6'b101010: cntr_next = '0;
    6'b101011: cntr_next = '0;
    6'b101100: cntr_next = '0;
    6'b101101: cntr_next = '0;
    6'b101110: cntr_next = cntr + 32'b1;
    6'b101111: cntr_next = cntr + 32'b1;
    6'b110000: cntr_next = '0;
    6'b110001: cntr_next = '0;
    6'b110010: cntr_next = cntr + 32'b1;
    6'b110011: cntr_next = cntr + 32'b1;
    6'b110100: cntr_next = '0;
    6'b110101: cntr_next = '0;
    6'b110110: cntr_next = cntr + 32'b1;
    6'b110111: cntr_next = cntr + 32'b1;
    6'b111000: cntr_next = '0;
    6'b111001: cntr_next = '0;
    6'b111010: cntr_next = cntr + 32'b1;
    6'b111011: cntr_next = cntr + 32'b1;
    6'b111100: cntr_next = '0;
    6'b111101: cntr_next = '0; // reset
    6'b111110: cntr_next = cntr + 32'b1;
    6'b111111: cntr_next = '0; // reset
  endcase
end

always_ff @(posedge clk_i) begin
  if(rst_i) begin
    cntr <= 32'd0;
  end else begin
    cntr <= cntr_next;
  end
end

always_ff @(posedge clk_i) begin
  if(rst_i | soft_reset) begin
    led_val <= 16'd0;
  end
  else if(req_i & write_enable_i & (addr_i == 32'd0) & (write_data_i[31:16] == 16'd0)) begin
    led_val <= write_data_i[15:0];
  end
  else begin
    led_val <= led_val;
  end
end

always_ff @(posedge clk_i) begin
  if(rst_i | soft_reset) begin
    read_data_o <= 32'd0;
  end
  else if(!req_i | write_enable_i) begin
    read_data_o <= read_data_o;
  end
  else begin
    case(addr_i)
      32'd0: read_data_o <= {16'd0,led_val};
      32'd4: read_data_o <= {31'd0,led_mode};
      default: read_data_o <= read_data_o;
    endcase
  end
end

endmodule
