`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: MIET
// Engineer: Nikita Bulavin
// 
// Create Date:    
// Design Name: 
// Module Name:    tb_miriscv_alu
// Project Name:   RISCV_practicum
// Target Devices: Nexys A7-100T
// Tool Versions: 
// Description: tb for miriscv alu
// 
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module tb_miriscv_alu();

import alu_opcodes_pkg::*;

parameter TEST_VALUES     = 10000;
parameter TIME_OPERATION  = 100;


wire [4:0]  operator_i;
wire [31:0] operand_a_i;
wire [31:0] operand_b_i;

wire [31:0] result_o;
wire        comparison_result_o;

alu_riscv DUT
(
  .alu_op_i (operator_i   ),
  .a_i      (operand_a_i  ),
  .b_i      (operand_b_i  ),

  .result_o (result_o     ),
  .flag_o   (comparison_result_o)
);

integer     i, err_count = 0;
reg [8*9:1] operator_type;
reg [103*10000:0] line_dump;
wire [31:0] result_dump;
wire        comparison_result_dump;

reg [102:0] running_line;

 assign operator_i             = running_line[102:97];
 assign operand_a_i            = running_line[96:65];
 assign operand_b_i            = running_line[64:33];
 assign comparison_result_dump = running_line[32];
 assign result_dump            = running_line[31:0];

initial
  begin
    $display( "\nStart test: \n\n==========================\nCLICK THE BUTTON 'Run All'\n==========================\n"); $stop();
    for ( i = 0; i < TEST_VALUES; i = i + 1 )
      begin
        running_line = line_dump[i*103+:103];
        #TIME_OPERATION;
        if( (result_dump !== result_o) || (comparison_result_dump !== comparison_result_o) ) begin
          $display("ERROR Operator: %s", operator_type, " operand_A: %h", operand_a_i, " operand_B: %h", operand_b_i, " your_Result: %h", result_o, " Result_dump: %h", result_dump, " your_Flag: %h", comparison_result_o, " Flag_dump: %h", comparison_result_dump);
          err_count = err_count + 1'b1;
        end
      end

    $display("Number of errors: %d", err_count);
    if( !err_count )  $display("\nALU SUCCESS!!!\n");
    $finish();
  end

always @(*) begin
 case(operator_i)
   ALU_ADD  : operator_type = "ALU_ADD  ";
   ALU_SUB  : operator_type = "ALU_SUB  ";
   ALU_XOR  : operator_type = "ALU_XOR  ";
   ALU_OR   : operator_type = "ALU_OR   ";
   ALU_AND  : operator_type = "ALU_AND  ";
   ALU_SRA  : operator_type = "ALU_SRA  ";
   ALU_SRL  : operator_type = "ALU_SRL  ";
   ALU_SLL  : operator_type = "ALU_SLL  ";
   ALU_LTS  : operator_type = "ALU_LTS  ";
   ALU_LTU  : operator_type = "ALU_LTU  ";
   ALU_GES  : operator_type = "ALU_GES  ";
   ALU_GEU  : operator_type = "ALU_GEU  ";
   ALU_EQ   : operator_type = "ALU_EQ   ";
   ALU_NE   : operator_type = "ALU_NE   ";
   ALU_SLTS : operator_type = "ALU_SLTS ";
   ALU_SLTU : operator_type = "ALU_SLTU ";
   default   : operator_type = "NOP      ";
 endcase
end

initial line_dump = {
103'h1e88592d984c690cac00000000,
103'h18f51e266e7dff015e00000000,
103'h22fd89520d06582ef800000000,
103'h0e6a324c64fb76556635192232,
103'h2eb6654386f8ffa77200000000,
103'h274f0147566331f3d600000000,
103'h0d659c4c851997375ebecfbfef,
103'h3e828f80ab68987eb400000000,
103'h149af90a36ce34cb3800000000,
103'h32ac623b3550c44be300000000,
103'h2620fd6008ebbd561800000000,
103'h1eaf2fbc3c981f914c00000000,
103'h00a5fa9722b91cf154af8bc43b,
103'h196afa3d42684cad9000000000,
103'h2480be2f430e4744b400000000,
103'h3a823f775d794181f700000000,
103'h0a1be050c0f9ffb13800000000,
103'h3e6e9e1b7a7c3f289400000000,
103'h3529a893c6981f795600000000,
103'h2ef2fa50c406bd94d000000000,
103'h03358d8fba30662896363ee800,
103'h1972207fe92360795c00000000,
103'h2a2af298ab58ee091600000000,
103'h017be42ac4cb0e88fe237959e1,
103'h1cd39351aef60121a800000000,
103'h325ba8a12e71e54c6d00000000,
103'h31071e6a0c45789e1a00000000,
103'h1a0b823bfea1213f4a002e08ef,
103'h06daf496f0a83fa95600000000,
103'h22a068138ab3c1e55400000000,
103'h2cd7c0dc908eb67c4400000000,
103'h02549243b22f1e8fce2490ec80,
103'h167284ea1f06df6c6000000000,
103'h1c38b739e05b71b01200000000,
103'h2ab2ab6ef8cdf69a3200000000,
103'h0abb56205406add412002ed588,
103'h1ef31f617eb959430a00000000,
103'h1131c80f0a74af635e5e8c55d6,
103'h22cbe26ca967cec4de00000000,
103'h2f33f364789996d3e800000000,
103'h0ca2b2305b65794090f3fdb86d,
103'h2acaca3f48996ca50800000000,
103'h136791b1963c1ed56200000000,
103'h226c27e8c106e914ac00000000,
103'h2b0a54f3d56e7ac64200000000,
103'h0e0dfb3f76daa2af0204511781,
103'h3aab0e3022e4f7a2d600000000,
103'h3c843ff630f2f2e24f00000000,
103'h3f645ad0ea9e01127100000000,
103'h16b2f071e7224108a000000000,
103'h24dc28c1e4869bd98a00000000,
103'h14ea58b4bb398c4b7000000000,
103'h34eb7b89de15b50d5400000000,
103'h3e8a9f7173000dc21000000000,
103'h2e4c0461a6eb894bee00000000,
103'h0294052b657628bd622b640000,
103'h1215924092c22d1f0800000000,
103'h02acd4631756324a6ec5800000,
103'h24442447a86bc48b0000000000,
103'h2cc6fd782a1898ee1600000000,
103'h1abfff660f5cbd35c05fffb307,
103'h1d7b2e72fc23baadea00000000,
103'h328c8fca56e3ba13fb00000000,
103'h3209b5acb35ee886f700000000,
103'h1e9f747d26eb78514c00000000,
103'h1891f08358f52dfe0000000000,
103'h0ea827377694a27b2640111993,
103'h1aa217ff8e2692fe7e00000000,
103'h1afaf14e9cceba35f60000000f,
103'h013f42eef870d23584d80a923e,
103'h0078c28d536bc38422f24308ba,
103'h3746e4a6d4ab06731a00000000,
103'h3b3b99bed423c9006c00000000,
103'h1cff090cca6aada74000000000,
103'h36334a9044a647661400000000,
103'h24d34f97e2a55072de00000000,
103'h241e5b1298d89b032400000000,
103'h3a8d2f8dbcabea9b0600000000,
103'h1966b1b022ca45ad9e00000000,
103'h3ce67b389d57753b5d00000000,
103'h020b9533f4be26eb7e00000000,
103'h23094a3272a4a2241a00000000,
103'h3eb2e9cbf4b037580f00000000,
103'h3c26cf1316b9818a8100000000,
103'h16f22995956c6b567600000000,
103'h247bab0390933a698c00000000,
103'h26a9ce95a68563ff2200000000,
103'h1c88297fcc010f02b200000000,
103'h292005f472aadd985a00000000,
103'h0b244dbf8f3307182600001244,
103'h3ebbcff437530d0c9800000000,
103'h18d8b62803775acc2600000000,
103'h3ef6ab5e80332ac05d00000000,
103'h16bf7e2d580be0e85e00000000,
103'h3cbb581456028c46de00000000,
103'h190a3f07ecc20a743600000000,
103'h38d080c7a87d62888c00000000,
103'h16c9ed47c087a1907800000000,
103'h0ecf3ab0385822582024110810,
103'h1ad7145f91220f9fe2000035c5,
103'h14a0f8831ef14a501a00000000,
103'h34e83f2f38c85eafaa00000000,
103'h16b7276bcc695732c800000000,
103'h32de3200835196620300000000,
103'h1c274c351808bdcdce00000000,
103'h2661b0b9cae6efce5000000000,
103'h296473ee290e3c036a00000000,
103'h36d08e554e6fecbd3400000000,
103'h088e3f1e76d460ab5c2d2fda95,
103'h3254adb56ca4ef00ab00000000,
103'h26020c1ab4332e1f2000000000,
103'h04bda6836687dbd48e00000000,
103'h2ee92da94e89e7ef4200000000,
103'h10e9157a93478e72aad0c383f4,
103'h1e8dec4c8130bc1bf800000000,
103'h2065f13d9119d1968a00000000,
103'h0ac5d2032ea7bde30a0317480c,
103'h02af9ab8110daf209c57020000,
103'h0ce0f1df9ad38123ca79f8ffed,
103'h194305231e831bdbda00000000,
103'h34bee9fd2b640dbb7600000000,
103'h3ee28cba42a712de9500000000,
103'h1a13de97f665fcdbbe00000000,
103'h1118b1997748899602e81401ba,
103'h24a0a076d05c682df800000000,
103'h228c9d0fa07519c76e00000000,
103'h251fac870415ba3e3e00000000,
103'h1e18b8da26a2574dde00000000,
103'h0d5a4ec34cc203d4e2ed27ebf7,
103'h0cf84cda6adabcaf0a7d7e7fb5,
103'h2a0b64b8f7350b725600000000,
103'h0e3436d5c32d584cc012082260,
103'h18ff60406e38bd05b600000000,
103'h2e8c8d7ffd6cf3db7a00000000,
103'h2ef4776e956c541be800000000,
103'h24916ccf82f8e19be400000000,
103'h1f5bba7d30ed590a7800000000,
103'h065ec530957ec5d9fa00000001,
103'h2acec3bf74da80572a00000000,
103'h22ab166a3a394587be00000000,
103'h1c804ab0e60809473200000000,
103'h0642d80208b31fb16e00000001,
103'h06842b2d27336a625400000001,
103'h389ffeaf6c7642645c00000000,
103'h26f517b972fa6d918200000000,
103'h3b523a0aac9a6c40f000000000,
103'h18627c0d528f83fa6200000000,
103'h1aa628724ee1be050e00a62872,
103'h0b60173ba7443a126200005805,
103'h2e14739680ea6284b000000000,
103'h3d633c324d4a79c05600000000,
103'h1f4188c87a5eed56d600000000,
103'h0e019363b6c229892200008091,
103'h2505d8115603b2519c00000000,
103'h3cf47f43a50545b55500000000,
103'h1f2da0364b0b1dc6aa00000000,
103'h3cc5ae7fc6ff9d0a4f00000000,
103'h101fe652642d3d4098f95488e6,
103'h3a7dd076a0f2ebc05e00000000,
103'h08e100503112d212c4f9e9217a,
103'h224f4df06a90a2896400000000,
103'h00bd389af571a2d996176dba45,
103'h0558608616c0f0ca0000000001,
103'h2ae67431967e2964f400000000,
103'h008759efdcd689eb0aaef1ed73,
103'h00b8e23786bcfe1ca2baf02a14,
103'h375c0d58c744580c7e00000000,
103'h00c0294406fd3a4404deb1c405,
103'h22a26e943d59479cca00000000,
103'h215b3dcf7e1970e0d000000000,
103'h24d10b2760bbdf750e00000000,
103'h2e8b308bc3171d448c00000000,
103'h0042903426e8286bec955c5009,
103'h0f533779567358f7ae29883883,
103'h1b7d4f9f56b5e92bd6fff7d4f9,
103'h0763473a650920a52c00000000,
103'h37605c19fe8670448200000000,
103'h0c45996584e9b77ee676dfbff3,
103'h389e2fa8bb4a1398e400000000,
103'h3aacaf17c68facfe6900000000,
103'h20c44f2bff2ddca72400000000,
103'h04625f84b8da8bbeea00000001,
103'h2cea275c589edaeaea00000000,
103'h10bc02ccdc013a6fa25d642e9d,
103'h3d1d8b3bcaeb61cbfc00000000,
103'h26acf051daa76498d800000000,
103'h0816e126d6c4efd4a26907793a,
103'h041face6bd71e0267e00000000,
103'h1f29b3164688c14d5400000000,
103'h001f1b11caa86e341263c4a2ee,
103'h3ebbe7a628d2214a5800000000,
103'h151da40f2af13c5c2200000000,
103'h26f1409ea8ad24024c00000000,
103'h3e4d9e7b7ccac8117600000000,
103'h20526a8c62bc08b01e00000000,
103'h2c2957e7a109a72b9c00000000,
103'h22f1819f025c11b7fe00000000,
103'h0266cf58ae85699fa0ac570000,
103'h1ea6e523d376eb3ea200000000,
103'h1ca3039f14ddba975000000000,
103'h3ca8c945f2849fbb2200000000,
103'h1e0aa0a4ce27a35a3600000000,
103'h30f1e1a34cd06ca02800000000,
103'h12500de06adb0d44f800000000,
103'h0a8bf4b4dacceee844117e969b,
103'h334c7b446e1cfcc8af00000000,
103'h2b34a52e38a8f17d8a00000000,
103'h2eed3bb82af56cc1f800000000,
103'h1e80df87172a11f03000000000,
103'h28e1723e44174da85a00000000,
103'h205f01be22982d2f7000000000,
103'h108582bb8b799f6db685f1a6ea,
103'h2aa1707aead8a12bd800000000,
103'h1ce7702a7b5e23e76400000000,
103'h1344bd8266ff94624e00000000,
103'h2b3a3809c2e7048cca00000000,
103'h0ea951fed52bc20f3014a00708,
103'h1ef10d1fbf65fa18f200000000,
103'h2896ec280f0f4c17c600000000,
103'h193c5f92ac0059378400000000,
103'h0ac8d78a1497455f92003235e2,
103'h10811190acd3a4f23ed6b64f37,
103'h149f45b0369c7c7c5200000000,
103'h28ccc5e7861d8e0cfe00000000,
103'h26fa9f565abcd3bd3400000000,
103'h3abfbe24c28999a4bb00000000,
103'h395881e56a8438fb1700000000,
103'h2e8dc2226443f71fd800000000,
103'h28e0906c5c9c79054200000000,
103'h3ef032738a2a3b27a700000000,
103'h18896e1f750acb940400000000,
103'h1aa6e2c672fafe078e00a6e2c6,
103'h02084e8d4a846c2702084e8d4a,
103'h07063359672b4eed7600000001,
103'h152e534d28339d7ac000000000,
103'h19613ed4ee39d0d42600000000,
103'h0e8f2864426824214e04101021,
103'h0e417e1a9ac962f63c20b1090c,
103'h361f22be69588b5a8000000000,
103'h053064dcf89a09751a00000001,
103'h037b77cfaeb92c3384f6ef9f5c,
103'h022eaee3b2e991107c40000000,
103'h1cab48edf56508e02a00000000,
103'h20806e52b693b7c3dc00000000,
103'h1cef9d2c953f00b1d200000000,
103'h0617f839f4bf6f048800000001,
103'h2529e457d2af0c311c00000000,
103'h36a0d955d8c7046b1200000000,
103'h3eab8617bcf0e8c2e400000000,
103'h1cf5338b7291c218bc00000000,
103'h2efe5003b33d48307a00000000,
103'h12b678ad0e327bbbec00000000,
103'h0f35a5c17c30cbbf9e1840c08e,
103'h08a5bb98cee7446cac217ffa31,
103'h36a79388dc1cea2e2800000000,
103'h14e6b3a966c2a5c6f600000000,
103'h03584f85dd6a394fd49f0bb800,
103'h2afab721f150ecf93a00000000,
103'h2284632ab2a93c7f1600000000,
103'h372af9619ea3f3a10600000000,
103'h3094355f812856cbba00000000,
103'h0767aaad3753502d5800000000,
103'h0c8c0cf426e7858cd877c6fe7f,
103'h0759abba2d4f303a0e00000000,
103'h1ecb3e2138db3d2e3400000000,
103'h376527540134e8e86000000000,
103'h045260b41e0027099800000000,
103'h39271fa116654e5d9900000000,
103'h184b0ec81ab7af11b800000000,
103'h334a3b1d54deceb2cf00000000,
103'h0a7e505aec29dd7ae8000003f2,
103'h02b28ca21e7418983cc0000000,
103'h114c1746eaf268f32a2cd729e0,
103'h3a9d50fd6ca4f5954800000000,
103'h36cd5966bef10cdc3200000000,
103'h21273f4af88e5dd9a000000000,
103'h2af53dc76f5bb7405e00000000,
103'h1cb5a5371082f68b5600000000,
103'h3d1b023bfa783452c400000000,
103'h1a716c1d162dd989d4000e2d83,
103'h315633d7d448dbc5ce00000000,
103'h3696b2d2eeba47e2e600000000,
103'h0b5a285961107bbaba00000005,
103'h1a95d23296a72e8da8000004ae,
103'h00ff5595a00156e70880563e54,
103'h3ab1b4be7a9729199f00000000,
103'h221e5bca3a967eaf4000000000,
103'h2c9b7e90b448336dba00000000,
103'h0abfcfe4d9668f37f60000000b,
103'h0ae5782004020dc8aa00000395,
103'h06a24974cec1ddad8200000001,
103'h3cf59978daa755cd8600000000,
103'h26911ceaa1499f425600000000,
103'h2a932f945d3f38bb3000000000,
103'h30975006c2d055a5d000000000,
103'h065d4e26ad63853a2c00000001,
103'h36caa2141efad540ee00000000,
103'h06819543e55823679c00000001,
103'h3377c12edd22c57bbb00000000,
103'h223e42bfa2a45abf9e00000000,
103'h3f68498a961c1bee7b00000000,
103'h388d2596795a5eae1e00000000,
103'h170a2509f6c2a838b400000000,
103'h12a9e9f92f4fcdcf2c00000000,
103'h30ee09a80559f2d92200000000,
103'h244e45455703dcd25000000000,
103'h1008df90c6f1e67a548b7c8b39,
103'h32862214eb402bbfad00000000,
103'h025332683a490b50723a000000,
103'h167a3594accf2d655e00000000,
103'h02a515936e225fcd98ac9b7000,
103'h36c1dc0c869c95624600000000,
103'h141ece454841aaf5b400000000,
103'h2cc4cbce7e0387023a00000000,
103'h3239f6bd132255478500000000,
103'h28d1817940e721160200000000,
103'h2205a197b32117d31600000000,
103'h267b6cabdaf2994c5600000000,
103'h2af4bec23ef83ae40800000000,
103'h009066202573a78fe40206d804,
103'h16132e940f6866522200000000,
103'h1eb70edb0ef8cc724600000000,
103'h024d886e650bfb065621b99000,
103'h24dc3ce5c4c309e16400000000,
103'h2cde98ed0710924fca00000000,
103'h03495b466ceccf358e56d19b00,
103'h26acea1218cb68229400000000,
103'h311c73e41a14c3690000000000,
103'h3e4f079780c1ad7b1800000000,
103'h14922d9ab2de215f3200000000,
103'h14c222d3712d28f6b400000000,
103'h2ebd802ec4bf56916600000000,
103'h20cda0f31a817964d600000000,
103'h149f6f32893ef9939c00000000,
103'h3a4f5ed1290c9a86b700000000,
103'h132c77667eac09b93e00000000,
103'h2ec8e68d38fb688a6600000000,
103'h24e6cf18ca27dff0e400000000,
103'h2243b137f8f0c67e1e00000000,
103'h08ad2ddddcd79596e83d5c259a,
103'h2ec2b43cff1b46cee200000000,
103'h0cd3a32688c874acbe6dfbd75f,
103'h350c7200f68b28e9be00000000,
103'h17360759835ecc104600000000,
103'h16373248f76b3e113c00000000,
103'h1553a4074ea1456abe00000000,
103'h1b388a7264d877b3b4ffffffe7,
103'h16a899c7382c1bbb0200000000,
103'h1577752c5264a62d6600000000,
103'h08b18ea2a80d3ff49e5e58ab1b,
103'h0c8ced83bc84b520f0467ed1fe,
103'h3240c418843643c39900000000,
103'h1220b66850c331475400000000,
103'h03654ee58503f55fdaee584000,
103'h1cb727575624abc82a00000000,
103'h308db4ea1889faadae00000000,
103'h0a9a864074412205041350c80e,
103'h376a88de26ced6ef1e00000000,
103'h243e80dbb0695d2f9200000000,
103'h2a3724a166d3e60db800000000,
103'h08b9c314cd1266e96ad5d2fed3,
103'h1b7d838d36498b8ad0ffbec1c6,
103'h15101af4be034e9f9c00000000,
103'h3e0c0f8bd880d22cd200000000,
103'h0edbea30ac90ed219048741040,
103'h2cbe2bbeea9cfcad6a00000000,
103'h3ee9f8d7fa78e6de1700000000,
103'h11191490a737129d02f100f9d2,
103'h3ac9027625210b74fd00000000,
103'h1009dd7d353a2005a267debbc9,
103'h12e7b531ae03227bc600000000,
103'h0f3e73c4410cfff8fc8639e020,
103'h30cc44f3d2f4b52aaa00000000,
103'h397b2198623328eeeb00000000,
103'h34641e4292ff6de2be00000000,
103'h1e503d688b7a8f7b2000000000,
103'h0a495c877edeadbdb200000012,
103'h093730d11f2eeb263e0cedfb90,
103'h29582e09a87847adbc00000000,
103'h1b789924f0af787edafffde264,
103'h191393bb5807a6888200000000,
103'h168d3c0f72803fad7200000000,
103'h3135cf89cc93d368ca00000000,
103'h3556aab1e3210f783e00000000,
103'h2626fe58d356df020a00000000,
103'h32fef88846ad89b3ed00000000,
103'h315732652ed4880cbe00000000,
103'h3b433faae0d380950600000000,
103'h27505c68d12ab2fa3400000000,
103'h24b45828cb6df2a51400000000,
103'h2ac5dd9cb0be4f0de400000000,
103'h1eabeb1d5572a736ae00000000,
103'h33657933013884d35f00000000,
103'h1649ba42dee46ff0b200000000,
103'h049bedf7d249e923b200000000,
103'h22ac70baa893a3669200000000,
103'h172f9ab42f2f915e6400000000,
103'h08eb498110dc02190c1ba5cc0e,
103'h1a8b683ea60b9ccd3a00000002,
103'h3f75701ff0f6e64e4d00000000,
103'h0cf31b67ca824e8cf279aff7fd,
103'h06a0580e0af7beace200000001,
103'h132996cd56eada14ae00000000,
103'h06be7259dc8b3222b800000000,
103'h294a3434b0b4c8f00e00000000,
103'h1758449c76733b49ea00000000,
103'h0e5e13b11ebd6f7e9a0e01980d,
103'h1d4ebcda7615b41b1000000000,
103'h08ca98268573c7cc30dcaff55a,
103'h22fb3c62a2c284a6a600000000,
103'h349f1be8aa8d1ccd2a00000000,
103'h24006aed4c88592fcc00000000,
103'h0a776e0d002775187600000007,
103'h346238f8e527e005c400000000,
103'h020f888b6e9f4e12c41f1116dc,
103'h3949f4eb2501870baa00000000,
103'h3d0cba7aa6110f971800000000,
103'h02f6f5229e5b04823cc0000000,
103'h2d090fd05c67befce200000000,
103'h04ba7890df5eb41f8200000000,
103'h036d685d0b67c3efde17428000,
103'h243167c04f223c80bc00000000,
103'h26506ba5d08fa4ddc600000000,
103'h04d72e8836c10c9e1400000000,
103'h00bca58a1d117843e6e70ee701,
103'h0709e07be2e8a6cc1c00000000,
103'h1c7957ee62a54c563800000000,
103'h0378743eaaaf2cd21a43eaa000,
103'h1f389d2d072884c07e00000000,
103'h170a3e5f48a0f8ff2800000000,
103'h32c4865da6d9962c2f00000000,
103'h30241ab23ce3d48b7600000000,
103'h1832dbd8eea85ae91c00000000,
103'h066a21c01ecc759b5800000001,
103'h3c4260a676ff51744900000000,
103'h18f435b8fc6973346600000000,
103'h3089df56f8abd3dade00000000,
103'h38c7e3de10a00993da00000000,
103'h20d25e008329e8ead400000000,
103'h3edc29973af1ccc8e400000000,
103'h184f68625ac42ac96600000000,
103'h2c6e7b0858a05460a200000000,
103'h132d974232efbcc2fc00000000,
103'h38169c66df5e37cb5600000000,
103'h1af16e54708bcf0d88078b72a3,
103'h18906b0b6aa26b746600000000,
103'h2ecfbc230493d9c8d800000000,
103'h36fec9fd9d2444d44200000000,
103'h1c8c0fa38af400f74600000000,
103'h34a5245700f2caf4e400000000,
103'h3760a47ede7eda986e00000000,
103'h3eaffe6f9323feef7000000000,
103'h23239d348a84a36e4e00000000,
103'h108b3cf0c834a1dde02b4d8974,
103'h00e5a7a1ea583f126a9ef35a2a,
103'h0ebeeceb7ae37c033251360199,
103'h30bc31247cc923a51c00000000,
103'h1a3e18cbca881090980001f0c6,
103'h0ef4a250fb4441b51422000808,
103'h2b036ae896825a80de00000000,
103'h02f5af836576fcd1daf8364000,
103'h16b117c34f7a67ba7000000000,
103'h36f49093d370173dd400000000,
103'h107c4b1968212f01222d8e0c23,
103'h0086601fde15bf94f44e0fda69,
103'h140771f82e920aae5e00000000,
103'h3602eb8aee186ace3c00000000,
103'h2c6e7c5b831fdcc66c00000000,
103'h0afb3c2d3a22c8515a0003ecf0,
103'h069dbb93e69144acde00000000,
103'h32d245a8f08c80da1900000000,
103'h0e1f3a8c372a3c6dfe051c061b,
103'h2c8c0c35eafc8216ee00000000,
103'h051ba630f81bbca32400000001,
103'h033c84d8e4a7c8d90e21363900,
103'h30e9e45ae8c36f0a0600000000,
103'h14c1804aeafff3e2ea00000000,
103'h24959e51dae9d83dd200000000,
103'h2a8578fbeeab5888bc00000000,
103'h161d1c7f1240f6da9600000000,
103'h29782f0c3ec66fd68600000000,
103'h26d3357c54e38c559800000000,
103'h3c18142a3c5bbb61d700000000,
103'h02084b60e22ef0de2a0e200000,
103'h1d397972214705086800000000,
103'h32311759e24f50694b00000000,
103'h1e0c41973e88c9db6a00000000,
103'h0743273672b9e1354e00000000,
103'h10a8fdb3d0c622cc8cf16d73a2,
103'h3d55d93996094a02fe00000000,
103'h0a520528a6b247b6ce00520528,
103'h16d6faf3220820f06400000000,
103'h1615d1f2ed5a26190c00000000,
103'h251acbbf4431210c2e00000000,
103'h0b290f8e9b46f2ff1c0002521f,
103'h16e99b14bf61bebe6000000000,
103'h04b2478b488ace4cfa00000000,
103'h20d51a1ade746961b800000000,
103'h01290db6a526b0ed0227df51d3,
103'h3ac3f45184fbcb07e000000000,
103'h34c099aac624d8be8400000000,
103'h36480d5100e8cd100a00000000,
103'h1643ea58f4a966bad000000000,
103'h1c66784deaf1740bd000000000,
103'h2684d14ac3355e64c600000000,
103'h36c803061e9bd6b2b000000000,
103'h06f401d18420a7fd7200000000,
103'h0cc96757bae8ab039074f7abdd,
103'h3e9040e9c0dcacd51400000000,
103'h308c78e08ea6142cce00000000,
103'h0324878a0d3655169043c50600,
103'h16dd3e30fcc2cdf71e00000000,
103'h267e9fdb7ee755812a00000000,
103'h36fcae5b16c493b22600000000,
103'h1520d1077d43338da600000000,
103'h3f7b48ca733fe1e8bd00000000,
103'h24988e848760b2f03800000000,
103'h0a9d29bfc4dbfbbaaa00000274,
103'h066658ad29748a3f3000000001,
103'h3f72bb283511b3fef500000000,
103'h28beff8bfa780cac1c00000000,
103'h196bf6dffaeac7d45000000000,
103'h0cf4e9eea2a9c7604c7ef7f777,
103'h2af2673c7d15be404600000000,
103'h3a019889480aa82ee800000000,
103'h0688d68232fd0f6b6400000001,
103'h0cfadc4f6efea7f4ae7f7ffff7,
103'h3616a97cf4877e76e000000000,
103'h1b4834eac2825ac64eff4834ea,
103'h0884688778990443440eb6621e,
103'h2abdab8f92e1392e0600000000,
103'h38f5968c5d65a1b57e00000000,
103'h3cb5000006234d451000000000,
103'h02f6c439fe18e3d16c3fc00000,
103'h00d18cb73ccde3d172cfb84457,
103'h128d8e627ec4a80b7200000000,
103'h3eaf31c3409634c2af00000000,
103'h32f422691223c3252d00000000,
103'h2451f6e050d2f4e86c00000000,
103'h127daf2902c717517e00000000,
103'h3e6e0f7d27190e31d000000000,
103'h2cf4a493f896bd5ad200000000,
103'h2a9efccff904ccd7fa00000000,
103'h3b1c49f464f9716bf200000000,
103'h0e60ae6a4e986e3bea00171525,
103'h08be21120ab4b8304e054c9122,
103'h3ab251149915669a9f00000000,
103'h26ab4def20d387aca800000000,
103'h349dbc359a85d8c14000000000,
103'h122898b8013126b06000000000,
103'h3b682d6ab6cee2e5fa00000000,
103'h3abd28b808f77b9dfc00000000,
103'h1ae5abb2055fa908b200000039,
103'h1694076d3e1cd1c0ba00000000,
103'h137389d8da027d72be00000000,
103'h0521ef2a709684dffe00000001,
103'h3ec7d01a030a0eb8d800000000,
103'h3ecd5a12472bfde34800000000,
103'h3cefb5cb44f3cdfd4b00000000,
103'h14148ef702c1280f9000000000,
103'h1ccfed02beb0dddad400000000,
103'h269559c752c56cd1d800000000,
103'h3686c46f2e9559d49600000000,
103'h0a6bfd14552ab39bea000001af,
103'h22125dc90ab1780b1800000000,
103'h3b699c58971d751f6f00000000,
103'h248647b9f82fd2e87800000000,
103'h3c384ceff2996f410f00000000,
103'h2a1505c1d71fb6fb0800000000,
103'h24a3369ed45803eafa00000000,
103'h324edc9b3f6d09acd300000000,
103'h3a2a55802310404ba700000000,
103'h369f3da6165f1ce6e400000000,
103'h0833dcc710897267085d57500c,
103'h2e207fd30728b00d1e00000000,
103'h127a2c8bce5c8cd42e00000000,
103'h1ae419903d7d0ca7360000000e,
103'h38ad237b90f739330500000000,
103'h28ff9fcdeadb52c34200000000,
103'h1f7acc2d6488763ed200000000,
103'h235285610c88160cbc00000000,
103'h24a74b3bea02e23a2000000000,
103'h36f34a49cc55679b2c00000000,
103'h351a9c1af2fcb2d71600000000,
103'h14ca642ae8effd20e400000000,
103'h020242479d0a993bd6091e7000,
103'h193d029e72d4fd66be00000000,
103'h3ccd2a9074d73fae5d00000000,
103'h125a05598d14424cce00000000,
103'h12d6dd438ae16cdd4200000000,
103'h2e5e4e695c3b7236ce00000000,
103'h3cbabcf5ee124f7a5800000000,
103'h3eee6b30dd709de3b600000000,
103'h0c365bb8982b5ad9a41fadfcde,
103'h265fb91d9719c60a8200000000,
103'h1cc488b9645021c31a00000000,
103'h013ba7cf8aafdae0b2f5c1581e,
103'h032364c96774639a1693259800,
103'h1e367c9ce6b00b69a000000000,
103'h11635a7aead370330647f523f2,
103'h26e05a1c0809eccfec00000000,
103'h070d349dd86d474ad600000000,
103'h0cae72b9be4da166de77f9ffff,
103'h38ffbc3f445ad604b600000000,
103'h112475f7d00948be748d969cae,
103'h2e531c80480904fdb800000000,
103'h26ef0a53982d7af58800000000,
103'h1ad8998dc8809775d200362663,
103'h151cfeccae6fa1c96a00000000,
103'h1c6aacca08483b573200000000,
103'h2ec15fc51c653a23e000000000,
103'h1b458db5bacfe6edeafffffd16,
103'h0c4a531c289146b3066dabdf97,
103'h2ebeba4c02d6d468c000000000,
103'h197b5cd311212784ea00000000,
103'h1e9d397dfedfe1d0ec00000000,
103'h208efd16d65b3ea3fc00000000,
103'h0a120762b4f87821fa00000000,
103'h366be61754877538d000000000,
103'h34e6ec50de997c9b8600000000,
103'h2f41d45b560562b2da00000000,
103'h00f7fb09caec4f03baf22506c2,
103'h06a699da392e235f1000000001,
103'h20dcade379261e68da00000000,
103'h1aac3e883eccb84312002b0fa2,
103'h2a8131dfe0a966268c00000000,
103'h0442743b3a55a4aeca00000001,
103'h1931d9f5a6d6d68eaa00000000,
103'h24475e18eb194ac9e600000000,
103'h2e299a7f434b24bf8c00000000,
103'h1ab53d0c269282d8760000000b,
103'h00968447d6bc1d57baa950cfc8,
103'h0d4ea21230715a63e0bffd39f8,
103'h03200aa67007deabb6c0000000,
103'h3d3c97fa3c5680bde600000000,
103'h1eeba8267e768b645600000000,
103'h1556d5aa7cb3235e9200000000,
103'h3d335d925a9ecb851200000000,
103'h1217c425eef5a12f8e00000000,
103'h2652ab776b28fec1e800000000,
103'h39041e2d3e40c2e7d700000000,
103'h0768b441a4936e5f4200000000,
103'h2f6c15db1c978c8c8000000000,
103'h056518a4230040ce2400000000,
103'h06871a2f116c56a94000000001,
103'h06e9dea1d4d16f4d6200000000,
103'h2ae01173dd58897c7200000000,
103'h2a6dd0d26242681e4600000000,
103'h0cfbd0ff0e227992227dfcff97,
103'h3ef627d4f8904a648700000000,
103'h06c1edf8468c1b639400000000,
103'h28e63d98048243388c00000000,
103'h2e4cf5560a443130d200000000,
103'h02d626a6352a6ec8d83531a000,
103'h10efa25ae277641ee23c1f1e00,
103'h22953973264d8ac51600000000,
103'h3abd13c3f73d2d1ffb00000000,
103'h1e291f4598d266932000000000,
103'h34bf9990148f7a571600000000,
103'h2ecd77f972b8999cae00000000,
103'h0e28e127e678332cc214109261,
103'h24c177765645ab263400000000,
103'h142c7457e56e8c4e1c00000000,
103'h1726eb908b3003c47200000000,
103'h0cd9fc65de5c781c566efe3eef,
103'h28054067f48363ace000000000,
103'h1a762f90405d6012be00000000,
103'h3055ab06a962a07ab400000000,
103'h12652a4182d8d00af400000000,
103'h10d12198b52e7b119ed153438b,
103'h04c07c9cc693a5532000000000,
103'h3a0d37b39664c6ebd400000000,
103'h18bc93451c2543889a00000000,
103'h3944bee197327b3c3200000000,
103'h0efb658faeef0e814e75824087,
103'h2845b190e733cd62e400000000,
103'h1af4c47df52f32f292003d311f,
103'h28c91af39e74e4837800000000,
103'h0ccfeca57969a9016ef7f6d2bf,
103'h1ec5ccd8a332c3f50c00000000,
103'h18ef7a6eae02b09a8400000000,
103'h07485af74ec87d732600000000,
103'h1316200366b7f7e1d600000000,
103'h174d8e10ed0052d92400000000,
103'h3eb7c0137f1672dc8a00000000,
103'h1424a2b0956400ed7600000000,
103'h385a02c0d31bc100f400000000,
103'h02475ab2e64063b1883ad59730,
103'h3835057e1e9a66725d00000000,
103'h2c392325e0e1c1254200000000,
103'h34a141bb1916c6a36200000000,
103'h10252151444fe9c942ea9bc401,
103'h14e96498faf12b845c00000000,
103'h36480e530a164cd5a000000000,
103'h388879325effb16e9b00000000,
103'h14dfaab51547bfc1a600000000,
103'h3686c6010ed038f40400000000,
103'h101f0cd162afe3a91ab7949424,
103'h36cda0775936a9aa2800000000,
103'h3d7be58bea55b67b8a00000000,
103'h1671ea62212356f2e400000000,
103'h3e38282c5c9f3c7ece00000000,
103'h08ae499fb21126e0ee5fb7bfae,
103'h2c5b14bd31494f0d4c00000000,
103'h3b5d96563af798acfe00000000,
103'h2a836ee22752ad6a3000000000,
103'h374883ece2b043c06a00000000,
103'h351ebfd88c33b2a29000000000,
103'h253e4ad1827c368f7200000000,
103'h0e556e77769af667fe083333bb,
103'h20bf3f879cd941398000000000,
103'h12d954582b2eafb0f800000000,
103'h12271bcb4aedef389400000000,
103'h12f119cddec74390be00000000,
103'h0b560e3870ee5f5c0a055838e1,
103'h1e9443dc82df7929e800000000,
103'h1f0129318f3587625800000000,
103'h285bfdbf2cc9cb3eda00000000,
103'h107e15dd8acaf47068d990b691,
103'h288e8d57f326f22f9600000000,
103'h027e7dfc42a5080d20fe210000,
103'h2ca3f602eb3395651400000000,
103'h029339486eb2136156e521b800,
103'h234d70fe5b5609644200000000,
103'h372e9ae3dce942acb000000000,
103'h0eb4ccd67f36b3ab0a1a404105,
103'h116e942e37654e8ee604a2cfa8,
103'h00da6ee7441a1b65647a452654,
103'h0a9c53049488af939a0002714c,
103'h314779ce94631e7ade00000000,
103'h152954439eff717f7200000000,
103'h31707d478e46eb4e0600000000,
103'h0ed1c1b0e2703f91a42800c850,
103'h02bbb5add2e0bcd932d2000000,
103'h0908c825a2b27e8a16dd5b57da,
103'h2f554c1ce46e3437e800000000,
103'h20e8bb622c76fc5d8a00000000,
103'h36ec6a391acc487a6e00000000,
103'h20d0d5e93cb503dc9c00000000,
103'h2a67c02372a16e15b600000000,
103'h1a6cde95927243fef20000001b,
103'h36e8f9653eda04226600000000,
103'h2d315caf5846e2b7f800000000,
103'h212ec3d60e2fdc1d3600000000,
103'h06cd99127a6138cc8e00000000,
103'h3edeb24dda8ffca29d00000000,
103'h36c9cfaba15d95b51800000000,
103'h04fbcfc1603c4802f200000000,
103'h235dabf4570617ae9400000000,
103'h3a20c0f3db01e76ff500000000,
103'h2c73d295fd5f93644a00000000,
103'h002479ed3680545824526722ad,
103'h3511694764f426ee2200000000,
103'h3e0470502418a0db5800000000,
103'h24f95ec8da2a0a22bc00000000,
103'h064de0a5d92e7a72e200000001,
103'h1e22b6dafd27d93bbc00000000,
103'h1cebb3fe4275b9e19400000000,
103'h3ecd51fce29870bc9300000000,
103'h3ad8fa1e3e8424bad500000000,
103'h0f131cb27c5176b7b6088a591a,
103'h21751882762a70d5f400000000,
103'h364cce34043d8d887000000000,
103'h2cbcf4a226b2a60ae600000000,
103'h22b13fcb1cff743eec00000000,
103'h12f701abc8bc68e11200000000,
103'h3a6734626b6da8ac2f00000000,
103'h2714f4a17e64aa57f600000000,
103'h39755aeb78cbdeba6300000000,
103'h26d535745ee0d35be000000000,
103'h1cf178de57562e475800000000,
103'h3f7b64f47d2b63bbb700000000,
103'h1e69fb62991cdc9a0c00000000,
103'h3724708b1898418e8800000000,
103'h2cbfb90f76023cf12000000000,
103'h38b12fdb2e26ad7c3800000000,
103'h00ce0a629ae6668bb0da387725,
103'h2307c18414979666de00000000,
103'h1ad9ba341465a0c97800000006,
103'h0aadefd5366d624d8c015bdfaa,
103'h28a8d2f293471c81a200000000,
103'h228a1c9b9cf50c56d800000000,
103'h2f02fcab869ddf496a00000000,
103'h10e17d84e927fbe508dcc0cff0,
103'h2a2d60abd72af8908e00000000,
103'h14c06054690c76157600000000,
103'h1d486c53d239d6c14c00000000,
103'h2a6e579ca6fa3715b400000000,
103'h20bc3eca8442a3698600000000,
103'h2e351e88eeb0fb062e00000000,
103'h22ba745cd16d39d0b200000000,
103'h2b79a0f1fea25859a000000000,
103'h1833049ce05cccb67000000000,
103'h0a2f0bb14ad66da86e0000002f,
103'h2adc0dcbe30972455000000000,
103'h1cf649b72c387df69a00000000,
103'h0ab2ddfc19148bc27e00000000,
103'h1acc3ef7740ad579aa00000330,
103'h36bc0d9b3ebdb375c200000000,
103'h34b54e845a89f26d3600000000,
103'h1ee70d64114600087600000000,
103'h232d580644fb4e8cd000000000,
103'h187e782222e25bf0e000000000,
103'h0e8d4bb3c50fb3f7240681d982,
103'h1f2611b29e8e2c194600000000,
103'h3e04d7b9ed1b77cd0c00000000,
103'h22deec4e0d41897faa00000000,
103'h2a9b5cd30a4661399600000000,
103'h3767814f2e254d87a200000000,
103'h20c1d1e498c0aa5aae00000000,
103'h37379a470f282ba9dc00000000,
103'h1aeeec292ee9fd8e740000001d,
103'h08ec9f44e52197d582e68448b3,
103'h240f9fe83f1083feb000000000,
103'h18f34ae646fd23439400000000,
103'h1aff218e2b0cc32bd4001fe431,
103'h0af4f5c482000e121a0003d3d7,
103'h1e0c61d05cff2fa04600000000,
103'h323451dae6f42564c900000000,
103'h0f596529070087352680029083,
103'h148b3ba2f834d9100c00000000,
103'h1cbd202f068e3e391200000000,
103'h02ee345b5b1979dc0cc68b6b40,
103'h11136dec78d69a0b121e69f0b3,
103'h22392eb2bac4ce666e00000000,
103'h2e93c8890ad83c52e600000000,
103'h037ca0986e116b05a04c370000,
103'h307ef283dca5338eac00000000,
103'h1657de7a5f21d4271a00000000,
103'h36f598d74ea0c6aaf600000000,
103'h226b8f8724f8a5255600000000,
103'h3cf2f13c9cee3dfca400000000,
103'h341f8680bf59cd83ca00000000,
103'h0b6defebfd4cbec066000016de,
103'h2f5d2002306c45412400000000,
103'h3944f53dbada352d2100000000,
103'h1e1b0875e837552f5000000000,
103'h054ae931e27c4a6d0a00000001,
103'h24c788ae409752e2f400000000,
103'h36b06d6bc4e23c14d600000000,
103'h017387566aa9c4c3160ea60cc0,
103'h356df670615a322edc00000000,
103'h0ae4aff760cdb985460e4aff76,
103'h22f2bc61573baff5a600000000,
103'h3ee304e020205fed0700000000,
103'h047d122202131c4e5c00000000,
103'h2a715192c0f6212e7e00000000,
103'h30334a88c47333508000000000,
103'h0e30f3746ee484e34210403021,
103'h0d4efc4d2017cf6c06afffb693,
103'h0c8021742f48c2e076e471fa3f,
103'h0ea767c9ba97bf2d96439384c9,
103'h1641e16fc717e0a1c400000000,
103'h0cc0dff916bf486b7e7feffdbf,
103'h2357adee6c0129db4400000000,
103'h27373ec438c209d45a00000000,
103'h24ae8ec79a19b7c2c600000000,
103'h293dbf6cc050f686fe00000000,
103'h048c387d64ff854e9800000001,
103'h0adbdb694c3d44bb580006dedb,
103'h0aed882990c97d38bc00000001,
103'h2318ecac9ca558a20a00000000,
103'h3c9547b6a692e0cb9a00000000,
103'h3811280f48abcd783700000000,
103'h02ca4d234441152edca4688000,
103'h1f4cef6fff523d3e2600000000,
103'h1474ea5ec01c8a616a00000000,
103'h322fc6191e6979d16900000000,
103'h18966f4bb4de64302a00000000,
103'h033e2dad260e2a4948f16d6930,
103'h2d38294cbea49994fc00000000,
103'h164eaf4dc0e2c7422200000000,
103'h1eceaf202c1af08ee000000000,
103'h1c2d1322c3699fdca200000000,
103'h3e99a16ea2384efccf00000000,
103'h20aac94f7f65621f9200000000,
103'h029eb8727cff038e34f8000000,
103'h10ad98245ca9ccddb201e5a355,
103'h222617b2de4885502e00000000,
103'h16d6e63e30f61d748c00000000,
103'h08ed16e9121c35276a7891e73c,
103'h39024b222af31b659b00000000,
103'h04c14c38f2e0324eae00000001,
103'h2ec8d29feae27d70d800000000,
103'h0ac6767b6ea3c9a9ca0319d9ed,
103'h38e04f7e5f6c9c49b600000000,
103'h10ed43e6e83312c5245d1890e2,
103'h1ada6a9e2013624382369aa788,
103'h10aa0ec63000a62a6a54b44de3,
103'h361d7c980adb10c88a00000000,
103'h38fd86b39c851f8eba00000000,
103'h2510a39452a29c26c600000000,
103'h2e3722b88aa022da6200000000,
103'h2a5e48072eb0c66eb400000000,
103'h31607e1e5ee7e9273e00000000,
103'h12e7d3c44946312e6e00000000,
103'h0711c590f8a6af4ccc00000000,
103'h04dbda380a8e83111400000000,
103'h3356b54dd0a048a20d00000000,
103'h3eb9798ad57c22da1600000000,
103'h13626ef648d2d827e600000000,
103'h1eb213ae868c51b2ba00000000,
103'h34903b77daeec0a90200000000,
103'h1a0eabe338a0d4578a003aaf8c,
103'h17093f28af310fcf6400000000,
103'h18d6aa96083fbbb29c00000000,
103'h223067b61e48fadb4a00000000,
103'h0778e57f391fa5715400000000,
103'h2462379fda500d277200000000,
103'h2f7c998fe2c8f2a6aa00000000,
103'h02d6b732872b2a46865adcca18,
103'h3679cfb074a7c3d66800000000,
103'h213c8d9fb97e7b08ee00000000,
103'h274f58b66ef84ab96200000000,
103'h0e2b1673ce34d8591a10082885,
103'h3d31fe77b684310f8800000000,
103'h20e0aa5204af47835800000000,
103'h3b0dd13542e145fb0e00000000,
103'h053342d1e2c1f04d1200000001,
103'h1c8d8cc79ccfc1825400000000,
103'h2a6c07cce00304543600000000,
103'h3cf9ca557c90911bd400000000,
103'h1268d2d926fc98e8b400000000,
103'h0899cba9e4f6633e3237d44beb,
103'h1c9a85fcf65f36175800000000,
103'h129e44a43ef901c13c00000000,
103'h053294675c9387be3200000001,
103'h1cc37d132f31cc627200000000,
103'h1b4ac8fd336460c9ceff4ac8fd,
103'h0c314afe8f27dddcfc9befff7f,
103'h3e10cec12972a6da2e00000000,
103'h0c83da41f6a3f1d8bc51fdecff,
103'h0828b22534b4c099e64e395e69,
103'h3731ead243389adbdc00000000,
103'h3463015c4a614d011000000000,
103'h1b06bec0829337d352ffc1afb0,
103'h374e6dfd76f6392f9e00000000,
103'h074addd450fcf7f02000000000,
103'h1b7fe887074b65ed96fff7fe88,
103'h3816403acc9643c1e700000000,
103'h183fcfc1e7162c48ec00000000,
103'h2e5f98789e2c6c83b800000000,
103'h147c591f776c3c45a000000000,
103'h00e47fb3e4cbd4be3ed82a3911,
103'h38e2ea0a39482dddb600000000,
103'h18f780a9782cad919a00000000,
103'h193883cc730f979bd400000000,
103'h0ee5c3350a0718454c02800284,
103'h285ed75be23f9c11be00000000,
103'h3c20196071255f46cb00000000,
103'h0b0e08f69a8436a2ac0000021c,
103'h080b902896a450031e57e015c4,
103'h12102f9fe0b258f9b800000000,
103'h01546b28eabde9224e092a259c,
103'h1ebe05f8bcce18c23000000000,
103'h16abd76b3d2283eb1a00000000,
103'h243df8e0dae089e3d600000000,
103'h14827350308c614f1400000000,
103'h2e84d6e1d6ca5a2fee00000000,
103'h06555335ab4ccd802000000001,
103'h1b4853749ad1a461f6fffffff4,
103'h091bdd976026f797a09e950060,
103'h297bc9093a6f4b0c3a00000000,
103'h1ea60eab028b28a39a00000000,
103'h011d21ccec06f1acd49209bce0,
103'h3a65d950caad0057d800000000,
103'h16d5886c4aca2224c400000000,
103'h2ab48294062ffb758e00000000,
103'h031ea55f5d0583e1da55f5c000,
103'h068fb9d786ba0675e000000001,
103'h16adcea78ad8abd53c00000000,
103'h3096059c506865acc200000000,
103'h10ae3806a61634544c4c01d92d,
103'h0ccbee52d6ac39f09e77fff96f,
103'h0ea3ab14e65a71f74401108a22,
103'h1c5413ac3326604a1c00000000,
103'h3b6ce1f042ca0b5f0200000000,
103'h3e9be4889f1e1f0b3600000000,
103'h1b772111988b00fb78fffffffb,
103'h1eaccf91d726e5841600000000,
103'h1508de5c329e0695ae00000000,
103'h0d2ef885904ad62784b77f53ca,
103'h237331ba2453b483b600000000,
103'h11426bea3082ad09465fdf7075,
103'h15388b9e52f5dec36a00000000,
103'h0cccb1e822384aad9a7e7df6dd,
103'h12abae597670d64bec00000000,
103'h3ede5f4e823d88340f00000000,
103'h1893bd4cd6e9368d8600000000,
103'h073efa0e94c795dc0800000000,
103'h1422817dec5b5328de00000000,
103'h1a76df39329a4d37720000001d,
103'h2508c52888bcceb56000000000,
103'h0283e1a56233adee92e1a56200,
103'h36c693fe463c73171a00000000,
103'h176499800ac054bc7e00000000,
103'h289cec394086e8bac400000000,
103'h04920da7d6eb823ace00000001,
103'h02badd04fe886e740eb7413f80,
103'h06201f79421a7c1be400000000,
103'h1645b6aa04d55920e400000000,
103'h24f236958cf5789a2600000000,
103'h0a8a38bbe33b2f442c00000114,
103'h2eaaa956472d65d9b800000000,
103'h14e5960c90b79e959a00000000,
103'h00f5dbe3be6247ebe0ac11e7cf,
103'h38fb9a551547ddf87200000000,
103'h123c880a943db9dc3000000000,
103'h34aadb99ce3954314400000000,
103'h26d0cdbea175dc3bda00000000,
103'h165907cf5520b7d5a800000000,
103'h1c291fd87af185944800000000,
103'h3736f1bdd34a8d639e00000000,
103'h1f7e17d46e73ad3c1800000000,
103'h273b1a26e4aa9ef9ea00000000,
103'h0518d44f0228b6ce5800000001,
103'h1ee8140b6863d0f53c00000000,
103'h0901e12b6e7ca5443ebea237a8,
103'h228f5b878d64b94fa800000000,
103'h1ec774dd95669a7b1600000000,
103'h1e284501f6f5f602a200000000,
103'h06ece61b96bd6ae03600000000,
103'h1d2e2c7974e5afe22e00000000,
103'h3ed42c26fad295fdc500000000,
103'h34e0c64f9700c2773800000000,
103'h22e3567ad4d4ee9e3200000000,
103'h26a3518648b5b4edc800000000,
103'h1f48fc73ec990b689c00000000,
103'h10c13d5f523c5ceee442703837,
103'h193a40c1f2855962d000000000,
103'h348832c2c34696c22400000000,
103'h1a8bd9b15c80d784160008bd9b,
103'h2a288c0890090a46d800000000,
103'h0e019b4eaa94e3f8340041a410,
103'h256003f796bd7000c600000000,
103'h3e050362a4bf0b4f7000000000,
103'h332ada51ca1f0f470700000000,
103'h3959bb87c92412a9ac00000000,
103'h2a1d80b5fb4eecfb7600000000,
103'h309eb5e4f4a8a8833e00000000,
103'h1cdef6635ec629393800000000,
103'h123e4628ce64df1e2c00000000,
103'h10c1a897ec43d5818a3ee98b31,
103'h0a93f8027e821baa5a00024fe0,
103'h370eeff05143c4424600000000,
103'h035011175ad7bc44c4a0222eb4,
103'h1cf6115c90e6ac351400000000,
103'h22dfe7235236bd4c6e00000000,
103'h264bd8946f2ccea90000000000,
103'h3cfb8e47d00cb5cc5200000000,
103'h2a83003ff9588e60c200000000,
103'h2af11e6d34541ca89200000000,
103'h3e95f9e6ded71ce88a00000000,
103'h0167a4098ac83b55be17efafa4,
103'h134603f8895e353c9e00000000,
103'h1f7cf24848c5d9462800000000,
103'h1c07fd409b0bdd3eb000000000,
103'h3a6a25217888cf86f800000000,
103'h229488581690ccc79200000000,
103'h121d20cb50faf1e90c00000000,
103'h0b6b9284b48f7a412200005ae4,
103'h1ec5e17cc6ac9b0c7200000000,
103'h2aa8fffbd2182d912600000000,
103'h0d1ceb4270de0f0deeef77a7ff,
103'h3e8bc8721a870f09c100000000,
103'h268a1fe2e6a3fa4c3000000000,
103'h14351260252fc2be4a00000000,
103'h14f8326e8ab9e2a13000000000,
103'h0499618adeeef5015400000001,
103'h0ec19fb0f2e7276fe060839070,
103'h3e8dd823368088fabf00000000,
103'h1289d353c54228abb200000000,
103'h323fb12582d000cee900000000,
103'h32e483f89759d422af00000000,
103'h24707e3b889985483000000000,
103'h0c7d01793a7e0940c63f84bcff,
103'h3acbad629eee877c5000000000,
103'h2cea5a1aec6b88f58a00000000,
103'h3262daf5e73736582b00000000,
103'h0274e119132190731684644800,
103'h0f04f07d06846b68fc02303402,
103'h3883875d48f94c821100000000,
103'h0e6da73316fe3cff163612198b,
103'h0a8efd610e81c45c5e00008efd,
103'h1ad1e4021cef6b8f760000000d,
103'h3099360c287e68f08400000000,
103'h1059d49843504cf2a284c3d2d0,
103'h0718b02374e982feca00000000,
103'h0b59500b044357970c02b2a016,
103'h2c895b820a5c07ba8000000000,
103'h3637cfe994b557c58400000000,
103'h05369143c23eb3478e00000001,
103'h041ed59cb97683312400000000,
103'h0a4a718cbcad1474e6000004a7,
103'h18d2153742cbea119e00000000,
103'h3d0f10a74d165b9e5d00000000,
103'h228abf5ee4e870d59e00000000,
103'h037cf147a2f7817cea7a200000,
103'h1e1c37a5448240dbce00000000,
103'h3c87681486ff32237100000000,
103'h2608f422251b69c8b600000000,
103'h3472f10560a2d1dd3c00000000,
103'h26d46f6586abc5ff6200000000,
103'h1cb82ea17c1eb704c200000000,
103'h189b2000e2f3266a4a00000000,
103'h3a997b28feab550bc600000000,
103'h3e3aa82e5746750ca800000000,
103'h08879b3312dff035a62c35835a,
103'h0ef3453c901a9863fc09001048,
103'h375215b058a233970e00000000,
103'h1d5c3b2fe69578d39e00000000,
103'h18acd5bc1ce78e83f600000000,
103'h28dd607df843c9b3dc00000000,
103'h062883a3d0f09f6ff800000001,
103'h3e15da60b8cdffedf000000000,
103'h1a98a9f140f68391c2262a7c50,
103'h15030805be0c5df27a00000000,
103'h04b12fce18a507e3ba00000000,
103'h064ff7066ca80fe97800000001,
103'h02bcbe2cb3593fb792be2cb200,
103'h3c2008e4b8a936bdff00000000,
103'h368fb18f3a65f4eab000000000,
103'h08a4621d7885fdcf6a10cfe909,
103'h076122952e15af5ea400000000,
103'h397722c476ba117c1d00000000,
103'h223659b1bc1b34114a00000000,
103'h065b8589b49256d5c000000001,
103'h2406af3116c8b0877e00000000,
103'h2ec788371e2436113200000000,
103'h314272b9432ae5424a00000000,
103'h2ed8914cb0f26d796800000000,
103'h200106b5e134e032aa00000000,
103'h2af22ca68e0d717f5a00000000,
103'h130788a8710e78353c00000000,
103'h3c47c9ec9a00a4dbca00000000,
103'h197a78aa2e082d843a00000000,
103'h14e2079a6b4ff770d600000000,
103'h1e57080a02ca701b0400000000,
103'h1ada80aed6ac77b56e000000da,
103'h315e9e2f77037fbf7200000000,
103'h34eae93450de006e4800000000,
103'h22c72baa003c9e9dbe00000000,
103'h156dde3ab42787d20e00000000,
103'h1ec10880d6eeb37c0e00000000,
103'h1d17b2866c5c91b6c200000000,
103'h2d4c5cfa4b1d9a379a00000000,
103'h3abda60be7354cbe0700000000,
103'h3e5676ef9281a9b85000000000,
103'h18ddfb4f4e3f4fc43600000000,
103'h1ec21165cc95c6b3ca00000000,
103'h2ec3c1b3e573c2031800000000,
103'h24fabec00335d368e400000000,
103'h2eb3658470f9951cc800000000,
103'h06ab5c0d14f453dcca00000001,
103'h2b39194984a7b9613a00000000,
103'h323a98890a53156e4f00000000,
103'h3d71eb31768c2eb7d200000000,
103'h36a2d2f6a8c6c740de00000000,
103'h06c80e98a738b2725400000001,
103'h1895039bdcdb8568fc00000000,
103'h36b50e0d62a39401a200000000,
103'h0b614736bd38979d80b0a39b5e,
103'h08d447a0f2eda5aae21cf10508,
103'h2b7ffa7d7e4eece19e00000000,
103'h2b0732c3072334829200000000,
103'h0e31ff0a30a32f001010978008,
103'h2c9562eedcaa61c31600000000,
103'h3ee66c7e6adc60cd4700000000,
103'h0e8662ef9671c3bc2200215601,
103'h25498de35658303a8c00000000,
103'h2cafe7d724de932a2400000000,
103'h0ec0a38e0b28210d7a00108605,
103'h1cadc01236d808e49e00000000,
103'h000ca0528498ac72a852a66296,
103'h3ac3b0cd60466c84df00000000,
103'h1859547261530cd76400000000,
103'h02171924da16bda4c42e3249b4,
103'h20ace6bbf57012172600000000,
103'h04db60c5b6872b3c0000000000,
103'h0a504754563411f7f40000000a,
103'h31183aba5c0f72bdaa00000000,
103'h30f6ebc5275fba120200000000,
103'h2745aee71777f4cc5e00000000,
103'h101b9d45076ee09184565e59c1,
103'h12259d9aecb48f789a00000000,
103'h313f10ae7ed02cbda000000000,
103'h34b83dd410f5ca588e00000000,
103'h0ea95fc60334db070c102d8300,
103'h3009624976ed18db1c00000000,
103'h3f1df445869678a11f00000000,
103'h0b02b2ff369fdaea9600102b2f,
103'h26dd3c1174bdcf301c00000000,
103'h06eca02abec0822f5200000000,
103'h1ce91d1f249dbe40c600000000,
103'h387c12b4aa8a5e6b8500000000,
103'h0aaee334c6737b8aa800000577,
103'h109f82e4feef8e3f54d7fa52d5,
103'h1450a4c4889e71741a00000000,
103'h3c9f84e4d93df4591b00000000,
103'h1078c370ac8e991da2f5152985,
103'h2cc57d872b2e1e027c00000000,
103'h0601c5dcfaa6e1732800000001,
103'h28dc7fa6e66c5efa5200000000,
103'h24f52dc9ed6e24d74e00000000,
103'h0e9c750a964aa47e340412050a,
103'h2071da4dbb3fd2482200000000,
103'h2eee210408dc4752b800000000,
103'h24d6c6b4aa4e21a07200000000,
103'h062d913c993c42a47c00000001,
103'h3ecf0042bd1309592600000000,
103'h30b0419102409a95be00000000,
103'h2c6dca32010f9ad87c00000000,
103'h1379747372bfdc697e00000000,
103'h12c161595f2da69b8000000000,
103'h0f1c579872a71b0ef202098439,
103'h0cb7e86d44687c68507ffe36aa,
103'h0d63141a9284d400c2f3ea0d69,
103'h3ece1c315e3cbc6e0700000000,
103'h1166cae3ac9fd08898637d2d8a,
103'h12a694a4eb6decb9f800000000,
103'h1a4edace7ad4b79da4000009db,
103'h337bf4f8ce7b4c428f00000000,
103'h2ae5cb9128ca27110a00000000,
103'h0eef72b21b461c09d82308000c,
103'h1f67068d072be79b0000000000,
103'h28b35205941b5a4d1a00000000,
103'h007ae9c0b28260da207ea54d69,
103'h000ca88cdb35b2dfb6a12db648,
103'h1ae48362dab09ca06800000724,
103'h3ce845d3dabd452d4400000000,
103'h33076291f6a1c8901f00000000,
103'h1aa8e02a328a0e63fa00000002,
103'h1e8010a2249170f5f000000000,
103'h3e07ddba7f3a51202200000000,
103'h394cf0001eba61c24700000000,
103'h2933cad5dcc23f7cc400000000,
103'h0aa4b40f940f2f7ce20000292d,
103'h10a70e3f3c42fa52be3209f63f,
103'h14e3b98f06e7ae625200000000,
103'h38dac6a1168ebca18e00000000,
103'h3694132fea7276309400000000,
103'h0a5c8f3ba24d3cd1aa00000172,
103'h1968059a1ae150019600000000,
103'h2f5b2a5ae43ddf3d3800000000,
103'h18dd0bbd3ca5e4d75200000000,
103'h2ed163502a010f323600000000,
103'h2912f7b4c4de1aef7400000000,
103'h3a35dc1af2af7e3f9e00000000,
103'h32969fbe5ac275f46300000000,
103'h269d483916f8520f5600000000,
103'h04a4ffe6088ef1cdb000000000,
103'h288ad2826e2c3a06c600000000,
103'h3e20235e72d139ecce00000000,
103'h2e77ea2eda5c0c6f3c00000000,
103'h36c8030e997c2fcdb000000000,
103'h04a70dbc08f419fc8a00000001,
103'h02b252703ebc1d0b24e07c0000,
103'h328ed11143632ac72d00000000,
103'h3cc75c2185157d376b00000000,
103'h207c16ff76a44e48ac00000000,
103'h0d24ebd9f56baa6a32b7f5fdfb,
103'h3689ddbf94e7c169a800000000,
103'h2551fa6c620cad439c00000000,
103'h162f945098968b033200000000,
103'h3eb17c7d7ce8856f9400000000,
103'h1c9f0f14921819c02c00000000,
103'h0f74631552c9963daa20010a81,
103'h23566459ae68a5523c00000000,
103'h0ecef0a13cdd08678e66001086,
103'h393002585e336cc13d00000000,
103'h36a92dcfac025d627800000000,
103'h04ebef84a6325fbad600000000,
103'h0297568bdcdb8d8a842ead17b8,
103'h3a1fc5faa0c77d0f2a00000000,
103'h12dba22aa35ed39b0600000000,
103'h1699dbbd1e7e9995a600000000,
103'h008a750a715a3bc04af258655d,
103'h07569be246f4177d6800000000,
103'h2cea3fc9477e8c87d800000000,
103'h36dcb74b4cd5286a1e00000000,
103'h1e4dc862f8bf68336400000000,
103'h3719153af09c1f7eb000000000,
103'h14d879904ee9e7e1a800000000,
103'h39166a6d8602fd1c9900000000,
103'h282983b4dadb76ace800000000,
103'h12fc052f94f1e11a6e00000000,
103'h2a6aa628fc1b64cf4800000000,
103'h12c32f040e1769fedc00000000,
103'h011eb4fbba821027dad06291ca,
103'h0a55b1a04c453f2be8000002ad,
103'h277e8f5f4e63f427a200000000,
103'h00c2d1ed98b9a5c7f0be3bdac4,
103'h2a1e7e7abf3835273e00000000,
103'h0cfc3b2fc0fb0714d67f9f9feb,
103'h3d1f3710aa19858f9400000000,
103'h3aa627193615c0bf5500000000,
103'h10e6bce9b434f7cffe58e28cdb,
103'h265f87e16edb1ee93600000000,
103'h3ad359ee00c1dbd2eb00000000,
103'h3b60b18a262163b45800000000,
103'h3003c9e5a0f4bda25800000000,
103'h1adbda111a556f2c7e00000000,
103'h328f0925cb5939122100000000,
103'h0c04140d643513233a1a8b97bf,
103'h0a9a82a958c41c490609a82a95,
103'h2b25aee7a4c830566a00000000,
103'h26064a526e62b2ffc200000000,
103'h2d401ecf5a8861e76600000000,
103'h16af066f808eac39d600000000,
103'h1ae20a58accecb093000000071,
103'h00dd3e98437dd178b02d880879,
103'h163b25d79d5fdbd15c00000000,
103'h07216efe5e3d1a699e00000000,
103'h3696645ef57840413c00000000,
103'h12da24c8bc99af3f9a00000000,
103'h329bb6ab3230139e8f00000000,
103'h2ebd245f060a38674a00000000,
103'h091bac7c78a5ef127edf21b703,
103'h16f274db276313718400000000,
103'h2362ec796f7ebfedfc00000000,
103'h200377b6457134c92200000000,
103'h24ae3b5a66d421429000000000,
103'h20feee1106d798f8d400000000,
103'h02b2b4392a85d4533c40000000,
103'h12e53a4f4a84c2644200000000,
103'h2688f52e8d37769d6e00000000,
103'h2200d1505e1cb0ecb800000000,
103'h2750466b06a5a61b4600000000,
103'h14258fd8e8a6776ba400000000,
103'h0c7f9bab0ef6bdd6aa7fdfffd7,
103'h12111e1aa31c4daf9400000000,
103'h38bf5176f09be95aa200000000,
103'h22132aee82ad07754600000000,
103'h360d7bd1bb6c58ec3600000000,
103'h1afe8a8b9e7f83dab800000007,
103'h200be6f5148cffac7400000000,
103'h16b52cb92e8b8a381200000000,
103'h0e0b79f28e97712d2601b89003,
103'h02ce2018254c9de65680609000,
103'h15104a18745817d8e400000000,
103'h3cdf73c5372637f10b00000000,
103'h133a27aa0d3682097e00000000,
103'h372c4cbc0815f5ceb400000000,
103'h016b0fb45a501d78c0dd96968d,
103'h3e01ea85907c6a34c800000000,
103'h34befd47d2e779e92200000000,
103'h34b2921390e9646eb400000000,
103'h3ebc1cae04a861b68700000000,
103'h2115c4c13a5af3ca1600000000,
103'h14ebd709391710781c00000000,
103'h1aa9633a592cd53956000a9633,
103'h335053da2f18ac428f00000000,
103'h0e9fa63088c20f7ce641031840,
103'h2449ec50fa1263571400000000,
103'h320b42e988b209879f00000000,
103'h18f96ebb6cfbf5d89800000000,
103'h2e0046cfdf0738c22200000000,
103'h0cc92e613800a77d8e64d7bedf,
103'h24a47949a700ee4d6e00000000,
103'h0731cdb9b2ca1caea600000000,
103'h16bb1802576e95f84c00000000,
103'h054b9b0d1ea063b1fe00000001,
103'h2adcc595745b7bb45400000000,
103'h376ede6b38a716c17200000000,
103'h34cb13efa283dc56e600000000,
103'h0895df6c58f2bac21e33b2d723,
103'h3d010e9b0cbdceb1c000000000,
103'h22c7b97e1453ae1e1800000000,
103'h02357b229054bcb92445200000,
103'h0327191df51c76373a40000000,
103'h1d0b71db7651f159ca00000000,
103'h00ad994ab8790a77be9351e13b,
103'h3aa36ed814847c533500000000,
103'h06ee011e9732159dee00000001,
103'h0455099c50d584760200000001,
103'h3a0e0373d6c385949800000000,
103'h294007c31d188f30ea00000000,
103'h2af68865962692a4c000000000,
103'h04df1ea5fe669a67dc00000000,
103'h2e9d395c685d22cd7200000000,
103'h2e1ed9a76c3c41737000000000,
103'h0cb909235ad97acfda7cbdf7ed,
103'h3f79cb440af854774700000000,
103'h30a127cc96b15d9aa200000000,
103'h0a25a722952b28deac0000004b,
103'h10e667ec04cc50ab420d0ba061,
103'h3280a3854ef1f7cdd700000000,
103'h1f133395e0d85fb9dc00000000,
103'h205721411259033f2a00000000,
103'h38c637caf26c36d50a00000000,
103'h14019f0012c358161e00000000,
103'h3e2efe030a898fe11000000000,
103'h0a34bcbfde8b2ee12200000d2f,
103'h28937ebbdeba2ce42e00000000,
103'h395e778ce8eee9a40d00000000,
103'h1aecc8741082685fea000003b3,
103'h0904a93c48e0dfecd2f23b684d,
103'h16a7b8e5a2cda860e200000000,
103'h0104f5732cd2519d2aeba3882b,
103'h15511ba4c37a0a82ce00000000,
103'h361faa36437efff5fa00000000,
103'h22cf18b496d01b9abc00000000,
103'h314c2f93ceefc5d0fe00000000,
103'h2a9b981030bede859600000000,
103'h27650b0f610b0e196400000000,
103'h24ad7e048aa6a6299400000000,
103'h3ac60c94710bb138f500000000,
103'h1ece60f554b92f3d7e00000000,
103'h329593dbd17f3bd1ef00000000,
103'h2667d4dbae4d9cc74200000000,
103'h24e0bc0522e330a31200000000,
103'h12655467894b057ec200000000,
103'h16a31c076f2bc183e400000000,
103'h28601f79409115eb6c00000000,
103'h2a6abfb2563431f2da00000000,
103'h0f58908e8094516c1c08080600,
103'h3c9166e96aff111e7300000000,
103'h16f5fec83a57a1acf200000000,
103'h32ebac9276e908965f00000000,
103'h26158c4f8cdf075e9800000000,
103'h18d3bd78c0cab3f10e00000000,
103'h3690ffc066e040409a00000000,
103'h0ea5e3b4feb3fdb95a50f0d82d,
103'h1ca3d03ff644fd79c000000000,
103'h3880c42984eae12ec100000000,
103'h13286c04228eb16eb600000000,
103'h14b0541f5a0f75983a00000000,
103'h14ec39f3ec37e19c5c00000000,
103'h0a6d1d4240e835bbb600000006,
103'h04d8e1bf54d46fafa400000000,
103'h22d357ab1e418cf1e400000000,
103'h18dd432f251a6eb13a00000000,
103'h3d1f104f86edc65c5800000000,
103'h2249132b9ecb098b7c00000000,
103'h1d4785b75cea19db0200000000,
103'h34878534ff332d06a200000000,
103'h32e1f363db7ab2bdff00000000,
103'h342a27ef0f0237f2fc00000000,
103'h163d6605c0e42b56d600000000,
103'h153abdf7760e5345e400000000,
103'h106b42efcd4bb94ba68fc4d213,
103'h27167aa6228677431c00000000,
103'h0cc3ea4f72f1ba32e879fd3ffd,
103'h3355854f9a0834d90b00000000,
103'h0ef57395a6cc1f287e62098013,
103'h36e11b275921a4781800000000,
103'h035339fc2717180dbe80000000,
103'h00b71303dcf8333516d7a31c79,
103'h182320e49f4b6d313c00000000,
103'h165b4dedde0280351800000000,
103'h2cb51f6f3725a119b800000000,
103'h282608fe4c80ef079600000000,
103'h008f25c279360e76cee29a1ca3,
103'h3843afb7e05c17751b00000000,
103'h10fab9e262eb3d379407be5567,
103'h1ed765269a2eecef7400000000,
103'h3834ff726a29a6d1d600000000,
103'h0cc8a83509010bf872e4d5febd,
103'h02b8686cc2360b6adc0d984000,
103'h189365dc0efeb39fe600000000,
103'h0a9d503ad0b71c0ca8000004ea,
103'h28d0e16b6a4a81e8b600000000,
103'h0e057e9474e7d2238802a90000,
103'h367027285cb8b38ef200000000,
103'h2cd9835c2abe32236600000000,
103'h34f9fb9ca12e594bc400000000,
103'h2764f5c5ce07dca7ee00000000,
103'h0eb7c2128301d8449000e00040,
103'h12c341ee2b66ce0a5e00000000,
103'h008cf3ed381e901ce055c2050c,
103'h1084ff380ae1d20b0ad1969680,
103'h2e84e72aca6ec5f84200000000,
103'h1086a7621cf3c5304cc97118e8,
103'h1aef35a3cb78ac5b18000779ad,
103'h1e7654025aff53bd3400000000,
103'h2adf446bf6ee8960fe00000000,
103'h02b6facdd564dd635aacdd4000,
103'h3682765fff4421cf5000000000,
103'h36c69e4d42fb1c9d2400000000,
103'h100a19f7b87d92fd22c6437d4b,
103'h203c1f032e44314a6400000000,
103'h04d30171ff4e4b421e00000000,
103'h26ae05b01e8a6a454c00000000,
103'h0c84268b635d6bb74ceeb7dfb7,
103'h2ad7da63ca0b71676a00000000,
103'h376fbf86968f97f2ce00000000,
103'h0355efeb81677256987f5c0000,
103'h2ec68a95b6d731dd2e00000000,
103'h3c9490f73b2d21c8af00000000,
103'h156e08c028f3ac5e6400000000,
103'h02d7187be4883d559e1ef90000,
103'h30a79a8e38f64615c600000000,
103'h154f4e7dbacd5e91aa00000000,
103'h35242435ea74f91fe200000000,
103'h3aeca64c7ec4479d9d00000000,
103'h263d65b8b2e86bd38600000000,
103'h08846b3aaed512200628bc8d54,
103'h2698cf4e541277d8b800000000,
103'h2c222c81dc96e3136600000000,
103'h326fd153022fb261bb00000000,
103'h2ca5e1f7b151dee39800000000,
103'h12b104bc62c1b0369a00000000,
103'h0ece9f59ce67922e4a23490425,
103'h26831d0aa31896eaae00000000,
103'h01674d1d30e736447c2741b0d6,
103'h0c9d5c13566a534f1e7fafafaf,
103'h3a951b4016d1a06c4e00000000,
103'h36f46c9b226efc7fa400000000,
103'h166c54e0dd0417bfbc00000000,
103'h24cb736b14f8845ade00000000,
103'h0a94e5446b64d93bbc00000001,
103'h062ff78a0f304ca6d000000001,
103'h243a064f58c531eb3a00000000,
103'h20482cd45ef529754800000000,
103'h314ed7b4452f2fc4a200000000,
103'h2aba5bcfe4775c990000000000,
103'h35562c9256c6344d4400000000,
103'h16b72f400080901d2a00000000,
103'h160d5b62f4d6bcaf8000000000,
103'h1c92b74a8a8debef8000000000,
103'h068f6fcb229b47527600000001,
103'h07525c98fe2dfe9d0000000000,
103'h0695d98404bd6e682200000001,
103'h3cb0131e8a0fcb012000000000,
103'h3e5838a890a5a4852400000000,
103'h209ba5850e55b7a3ae00000000,
103'h030d10fe8cadf04c4086887f46,
103'h263beae02d4995d14e00000000,
103'h167a8fc2ef56a6cfda00000000,
103'h175ed92ad69291b00600000000,
103'h2498da366d0d2172f600000000,
103'h3e80cb8e436bfa9dcc00000000,
103'h04b252b76704d4d43800000000,
103'h3b3a80b06485a0627a00000000,
103'h065540596937f319e000000001,
103'h3f7d2175657273ca4500000000,
103'h3810fd2f2ac7b423ad00000000,
103'h18a9adbd2a44d5991000000000,
103'h1cc7feada355d2c83c00000000,
103'h0b1e42b7fcff808566000011e4,
103'h1ae6fa8c98c77f33080737d464,
103'h16776684e2e5c1eb0400000000,
103'h3d4ca8163eccbc779e00000000,
103'h0677bc6fd44422fc8000000000,
103'h0aa2514ed290cb12be00000000,
103'h28946560d90887829400000000,
103'h2a6c3b5de2aad8d16600000000,
103'h2910cdd28d3f3e323e00000000,
103'h3cf98343b6ab79902000000000,
103'h227303c79ebc4762ac00000000,
103'h20f50bce1cb5caa66200000000,
103'h0221eca5ff28ce6e0221eca5fe,
103'h2e8e0bb0211dda3c1e00000000,
103'h12a5a44a623fc6e21c00000000,
103'h1479844750cdd2923c00000000,
103'h32032eeaa27376dc9f00000000,
103'h0eb5a7fbf6ecfb23f0525191f8,
103'h0c85fb4968f02a0e927afda7fd,
103'h2a961578f8a5d20a8a00000000,
103'h1b74023ac42bcd53f2ffffffdd,
103'h2ec565d92ec1e2ccea00000000,
103'h3903c49b8a35e507af00000000,
103'h2b324d6c78fb4ae0de00000000,
103'h1706a847f0ff0f7c6800000000,
103'h0406d0775b315ce8e000000000,
103'h22c8db73b1380530d000000000,
103'h0ac0cb77b63ed5a82a00000303,
103'h2ab4065c9907b11bdc00000000,
103'h3aa650bde4c87c939200000000,
103'h26c9f8080e7c82f02a00000000,
103'h0325a4830a22d3ae0e6920c280,
103'h14c026a630eccbb61e00000000,
103'h3f6259e5331270392900000000,
103'h0ecd09b7c6d296df5860004ba0,
103'h2cb43c7a8534f0c48a00000000,
103'h14be42eb5301fa7c5000000000,
103'h2cb515123eb636f6d400000000,
103'h36be5772537479e22800000000,
103'h069a30b1be298ef46600000000,
103'h1aaafab5b4e7e666ba00000002,
103'h02bdbf35fa82171878d0000000,
103'h2a86baad172d11ce2e00000000,
103'h24c4300658ead1042800000000,
103'h1c2b345402718bb13e00000000,
103'h0a7a1f086735bbb7980003d0f8,
103'h354b20d54460f00b9a00000000,
103'h324934704edb0f140300000000,
103'h0a32190f83262fe946032190f8,
103'h268c895ff66f64599400000000,
103'h281cb56800a17d691800000000,
103'h2e0dd17ba72e06c90e00000000,
103'h02d9fca34e4abc310e7f28d380,
103'h1acc57b43d588dacb60000000c,
103'h292e171ec0328a500400000000,
103'h383153f25afee2044300000000,
103'h2f62978f052cf9230200000000,
103'h32de975cbc5e4d155d00000000,
103'h34b324d72ac0e4a46000000000,
103'h36ba3ca19c9f7c011c00000000,
103'h14c036705252a0d84600000000,
103'h34f32962090cdd79e400000000,
103'h128469691ccd13ea3600000000,
103'h18d68e1492c03d4c3e00000000,
103'h3cc82ec12544a6b55d00000000,
103'h320c7045fd1b34c9ef00000000,
103'h335d8f44bae3638b1300000000,
103'h0e7bc22dacefd3d10e35e10086,
103'h3c5a3262de4d6315c800000000,
103'h0e7d494d6cc92543762480a0b2,
103'h1cbb9501e82357a65400000000,
103'h26dd444176a0a0f3c200000000,
103'h1ceec752145c35f5aa00000000,
103'h314dad787b397a372200000000,
103'h3375b8e2572841893700000000,
103'h1ec11bf28775ef01b000000000,
103'h00ad1ff67aeba7e406cc63ed40,
103'h36f559f018acc3d68c00000000,
103'h27770e20d859e3cd0600000000,
103'h2d2103dace4f3dbd1e00000000,
103'h3940e89674c64bddf700000000,
103'h014c753620e74fb8c419e27772,
103'h1e04c5ac5828384f3800000000,
103'h1616f9ef9874ad855800000000,
103'h1b786beff9797331b2ffffffde,
103'h14a029ce4e906d214a00000000,
103'h2caf37656808d9114200000000,
103'h1ee67d4bbca902df9000000000,
103'h2a9270b76b583a44fa00000000,
103'h2cb7d754c83eb790b600000000,
103'h3e6dab1372d128482000000000,
103'h392c57e36088ff9ceb00000000,
103'h2e940792def6aab05c00000000,
103'h1153f18756230293bc987779cd,
103'h3a52930c84b70a269a00000000,
103'h16225cd9d40afbadf000000000,
103'h147b26440f5d8eba7600000000,
103'h2eca9a5ea67feb944a00000000,
103'h213d110cfafb11d85a00000000,
103'h166691e1e8c5ac370000000000,
103'h209b0e64c902bd43fa00000000,
103'h3a2d19a21e694f25e200000000,
103'h3b3f1073c1045d8aad00000000,
103'h344c191dba31772cca00000000,
103'h191ecdfeb67087a08a00000000,
103'h04f44023aabca0be4600000000,
103'h0e33016e82db6ebcfc09801640,
103'h1a76204406cfaee0a600000762,
103'h20eab6465702b04f2a00000000,
103'h1ccfd3e93078d0933000000000,
103'h0371924a506386d986c6492940,
103'h2ceebf686c335ac2b600000000,
103'h1e3b9b672ea4ed0d0600000000,
103'h248b27b51c93ac757200000000,
103'h1d5384963acf47dca200000000,
103'h227f6850df5a6f91be00000000,
103'h16dea6ce3aadf427f800000000,
103'h38e2d2589e2d5c78d600000000,
103'h377aaa58750c03471200000000,
103'h2ee1ca34eceed59fb000000000,
103'h04a359a323697ff82400000000,
103'h1712dd39514b4a2d1000000000,
103'h06afbd4854eea3d03200000001,
103'h2b58a09e6d0181098200000000,
103'h3af0599432b13e51d700000000,
103'h2cf192821e09def04200000000,
103'h2e3e159d18fa38847600000000,
103'h07793c8846ebcb069400000000,
103'h08b5e47cf429e0a3ac4e026fac,
103'h3ea3cac37aa31d2bf300000000,
103'h129b8ffa455901a8e800000000,
103'h008d8db582fccc6c62c52d10f2,
103'h336b567756985c66a700000000,
103'h1b72ffdcd725ea1c2afffffdcb,
103'h3e1dc66e489140938000000000,
103'h25218ea8a50440705600000000,
103'h0f22234f622206de9e11012701,
103'h0ebb145cc643958742018a0221,
103'h2579ef865665b8d6a400000000,
103'h04ca0b436520cd336c00000000,
103'h071e6770ca9abcb9c200000000,
103'h2c94ca7cce64c7fd2600000000,
103'h184ec31014832f6df000000000,
103'h1a6e747a0017f9eabe00000000,
103'h00aef3175966bcfad40ad80916,
103'h328a2e6e72d53174d500000000,
103'h30ca31c2b484248c2e00000000,
103'h048d6484e60e52faa000000000,
103'h1a689131d6d884bd54000d1226,
103'h08aa7ad99c65e9423a67c9cdd3,
103'h28c195f636ce7a741200000000,
103'h3f5cd59eff78f54dae00000000,
103'h38066842673a8b43e400000000,
103'h0a887fa3249760e2e20000221f,
103'h397080461e9dc9254900000000,
103'h1c26fb5d292648c86e00000000,
103'h3f566bc1e296c90e8d00000000,
103'h08c0676a7ebdc46bb43ed180e5,
103'h36c1c3f5fe14302d9600000000,
103'h0360e9a6c6d4979816a69b1800,
103'h3726581ffc965b8e1400000000,
103'h0e828fa7bef74534da4102924d,
103'h249c8b9b351d9d54d600000000,
103'h38cab7bc42a02cfc9400000000,
103'h12cd7b75663cb897c800000000,
103'h28669abc9f0770540c00000000,
103'h3cf6ff38b0d4ebc97200000000,
103'h04a50109993b86861200000000,
103'h10f32fd7143285bec260550c29,
103'h057e173c5ad786c85c00000001,
103'h16106ef5aacab69f7000000000,
103'h1877b2786e48cddbca00000000,
103'h341a7c8145593cd17600000000,
103'h26efcc48ded0ef49e400000000,
103'h309ca2d8d2eb6bcb2a00000000,
103'h2614300838db38140800000000,
103'h0cd48b136a77daecda7bedfffd,
103'h36ee22f0108c0af51400000000,
103'h3ed8aa169d6096087e00000000,
103'h18ae9d08524eb8f88e00000000,
103'h2c5fc80e1127630f2c00000000,
103'h2a88ce00aad600177e00000000,
103'h3a3ddee85735c8259100000000,
103'h275385d882be96263a00000000,
103'h24b7e5c13cfc750e9000000000,
103'h3543a8b9224ffae71200000000,
103'h2ea56bc88607e0a84e00000000,
103'h013cf6fd7c4b896170c4402f76,
103'h12931858aaf0f529f800000000,
103'h22e5aec26b2dec277400000000,
103'h128840133ec104801e00000000,
103'h0b32b20c60a6b3428a04cac831,
103'h3e28ad66f32ef355c800000000,
103'h1f0f9deb7f61a5622800000000,
103'h28247a977c8a52c91a00000000,
103'h30fa5bc39a99f0b49800000000,
103'h1876f03242be6b4c1600000000,
103'h322277f6b2b8c70fb100000000,
103'h0c2fa51d4b2fb741f497dbaeff,
103'h22c7250cfe522f38a600000000,
103'h12f895b14a81d455f200000000,
103'h06e871a1ad48f962f000000001,
103'h2e9114a1bf418f143a00000000,
103'h21696ee3c72a00b5e600000000,
103'h1093f85e74bb1557a4ec718368,
103'h0b40562f1424843b6a00000501,
103'h3135ad62a4b87c99de00000000,
103'h156c93aa6ef8d2c8f200000000,
103'h00cd7aa81e2e802b967dfd69da,
103'h1ee976fd729b13d60400000000,
103'h1229f78e32688e7e2200000000,
103'h2922f4b8d352057b9600000000,
103'h2f14c4ac647bfd09c800000000,
103'h103514cb8c9ef1c29acb118479,
103'h26f078c0bab3b66efe00000000,
103'h31146b340ce8cb3a8c00000000,
103'h0a8a6322f2d943fb4608a6322f,
103'h0a7c581ba2edaf2f52001f1606,
103'h170d3ed6ef7812524600000000,
103'h1d51dc0138f46a6de800000000,
103'h317f44660e01a944d600000000,
103'h3685f0c62a5385460e00000000,
103'h1e7a4c559ad2c9ac1c00000000,
103'h36e6ba375158ba724800000000,
103'h05479286f0d306c7e200000001,
103'h22aa141b66b9c0ff3400000000,
103'h2a601af5eb0153862400000000,
103'h0ce8eb7c8cab67a18a75f7fec7,
103'h00ca7675760b8297746afc8675,
103'h257f083644f46e140200000000,
103'h2eed5af644bee4897800000000,
103'h255d013c6a3decbfbc00000000,
103'h26780f24192b47b60200000000,
103'h1e9e9fa33c8848f26c00000000,
103'h1cb99e36620058168400000000,
103'h1e938153029ef7b9c200000000,
103'h0aab512f5e5895f0240000156a,
103'h0eee68c1bcec17432676002092,
103'h10b9c946869768728411306a01,
103'h368581e1d485d1344000000000,
103'h1cf03236e63f9a7ac600000000,
103'h22b3787c1cc51c5c9c00000000,
103'h2262d60478b54e938200000000,
103'h2aa99bff5b68c70f9e00000000,
103'h0776332e7ecb9d141600000000,
103'h088264d86975391372fbaee58d,
103'h2753b2deeeeb6c41f000000000,
103'h3cda4f78f76dd11a5900000000,
103'h2ec9b3229cc183f94600000000,
103'h1e84b3e0589bd3723c00000000,
103'h36b4edb189658694d800000000,
103'h3cd093c4a6ea3a753100000000,
103'h395a0af21e9f2826b900000000,
103'h10a50618db6fbbeb609aa516bd,
103'h028bd4b1d4c9c6dd7e00000000,
103'h3ad829dfa46eccf65900000000,
103'h1a0eb982a6faa1a82c0000001d,
103'h18e4714c62d2cb87d200000000,
103'h3229e5017ce1850a7900000000,
103'h1f391f9416c5f656da00000000,
103'h30b7271d08efdb585800000000,
103'h2a2fd04e2728faec6e00000000,
103'h057b450718e022097600000001,
103'h1ca83eca820ff2579c00000000,
103'h0a9b2ee4c68b375eb400000013,
103'h017dfa576433762936d8b8404d,
103'h1e89c0b66ecea50dfe00000000,
103'h1375a91ef14c9f656200000000,
103'h0b7183df0ed6601bd000b8c1ef,
103'h08f895fde04c093ac05a4e6390,
103'h2ab31e45eabd8d19ce00000000,
103'h3a3c4b9bf2b62317b000000000,
103'h3c1218575c69415d9b00000000,
103'h0abe452e98a58cf98e00be452e,
103'h3ab67b4094b7a550ea00000000,
103'h166c3e6c5e75ea7f8200000000,
103'h24d824afda2c65c01600000000,
103'h0ead4c50f098a42c7644020038,
103'h132800eb9570c8dc5000000000,
103'h285a5ad7231e152d4000000000,
103'h1e029f4235461618d400000000,
103'h2ed7496d5ea070eff600000000,
103'h2e4497c4fca310322c00000000,
103'h0322aef8ed7a599f8a2aef8ec0,
103'h3a1edb5a1abef1648600000000,
103'h27611dd41ee1a05d7200000000,
103'h3143d13e19007bb78e00000000,
103'h36c994da3f61998bac00000000,
103'h2ac9b215eea56ac9c400000000,
103'h3888c0b6256effa40200000000,
103'h24296fb3cf38b1b9f000000000,
103'h28ca9a6906c172701400000000,
103'h2acd5ea9eaeae223e400000000,
103'h1a758db492b57c8cea000001d6,
103'h2e8cbc633c82db36d600000000,
103'h12dc9ccbd6f868eb6800000000,
103'h3eedefa48685254ea700000000,
103'h14ea24a11861c21a7c00000000,
103'h3c9bd62a964fb1bf0200000000,
103'h22d062eaeb39d6601c00000000,
103'h20fd5896a8d5ac8ab200000000,
103'h22af73910aa60f759e00000000,
103'h3ec350a5eaa3680c4700000000,
103'h3326df79ce52db9d5100000000,
103'h10c444adcd162c433cd70c3548,
103'h1637566c7f3d0bbd0a00000000,
103'h265077a0ce01506ad600000000,
103'h220d00e16538a6d75600000000,
103'h2d1c65bf4c891e782400000000,
103'h0441f6e06e961f598a00000001,
103'h1aa493be9cb28518d6000a493b,
103'h3f088107a0f47bf94500000000,
103'h08a51527fa990fb7e01e0d480d,
103'h1ecac7c078a190bf8000000000,
103'h248699b28246a5e77a00000000,
103'h04f4f0bd61116da7f400000000,
103'h0657c3c18498075a7600000001,
103'h0153a67d8a8cf817d6f04f4ab0,
103'h34f119f910e4bbd95c00000000,
103'h2ad5335c11386256e600000000,
103'h02caba6707297c4ff618000000,
103'h1e5848cc70feafac0600000000,
103'h0472cf49b2c96a130c00000001,
103'h3a7211a05121b2df7f00000000,
103'h00a9b64dd4948229309f1c3b82,
103'h0e0ad74b4f0693c9820149a481,
103'h0d6aa7f4d0b04a1756fd77fbeb,
103'h3c93e2b15ebb2162a700000000,
103'h3eded04d6b25c9577600000000,
103'h16be4012a6b9ac08d400000000,
103'h3ca443a166987c563e00000000,
103'h333a91477c56bc68e500000000,
103'h068c005038fb000a4a00000001,
103'h050338b06a359151c600000001,
103'h29341d1970c191a1fe00000000,
103'h34fd7dd8b4c4ca526800000000,
103'h3a1d9b00dcf8e76bd800000000,
103'h3a38b83350f665448c00000000,
103'h228966b78d1400456a00000000,
103'h3c9ba6ddc64cb878ba00000000,
103'h0872b15668d61f304652573317,
103'h3242a33ae471c60e0d00000000,
103'h2f08fa63eee477647600000000,
103'h34e351d260271a9f5a00000000,
103'h020a61b98e30150348530dcc70,
103'h390790d1051366d5ab00000000,
103'h137685f6861dc88f3800000000,
103'h1cc9f2807e2559603c00000000,
103'h064479a9d09bdf56c200000001,
103'h3eef15d66c65d1d74100000000,
103'h3cad18d8b2aa4b811200000000,
103'h3e88e46a329961577e00000000,
103'h008a095bef467a3032e841c610,
103'h12270da46ccf5e9a6400000000,
103'h1029e3c42d5967f652683de6ed,
103'h02d70564fe80759abe80000000,
103'h271d885d50aa595eec00000000,
103'h38aa8585d2815ec3ea00000000,
103'h3906e148ba9ee7213b00000000,
103'h24bca501f3496ca70e00000000,
103'h0ef2de55eb504defc8282622e4,
103'h0ad37108ce0cf2f1ba00000003,
103'h1935627f9effd147a600000000,
103'h21363b17a8d342507400000000,
103'h1a808056c008a4d01200202015,
103'h011b1385a03edfe7baacf9b6ad,
103'h36c299a63abf603e7a00000000,
103'h0969f10e7cda73c41ad9c16533,
103'h04e48ac7329d0d6a5600000000,
103'h3e67c94ffb06fe78d200000000,
103'h1a29e7c07eeb894004053cf80f,
103'h30ab666f7e53528ffe00000000,
103'h030758e2997d3a507e00000000,
103'h070058c00928a0bffc00000001,
103'h050057164b2ff9a29400000001,
103'h02ebdeac913052629cd5920000,
103'h3e2ab8d2d530a978e600000000,
103'h12e6cd49991c88257600000000,
103'h2ecb8280564740f84a00000000,
103'h14e03159aa2e0e41e200000000,
103'h0a25329598f990c23a00000000,
103'h169add4a6ed9c21be400000000,
103'h382d1024b8fef4b17d00000000,
103'h320683f74e99d1fbeb00000000,
103'h170e060bc8c6e220a400000000,
103'h140f18e27acd6617f200000000,
103'h3ee9edd512db6c23bb00000000,
103'h22c3b77926ea85063600000000,
103'h1637531924d472db4800000000,
103'h1171d0d9c8982a546e6cd342ad,
103'h0779b4b25ecf7d6d9200000000,
103'h0e5d04aeae414e475a20820305,
103'h3d2ad9b136bb02f9b800000000,
103'h10cd218f051807a868da8cf34e,
103'h2b0793c14342e1599e00000000,
103'h25118361121002e8a200000000,
103'h0c5cc1483c1796a9e42febf4fe,
103'h2a63022920291a0af600000000,
103'h0c814ab26c85db533442edf9be,
103'h32e2749556e8dd7c5500000000,
103'h2953a160e56a282ec200000000,
103'h1cdc64d6564c9cc41800000000,
103'h328e4256bea03e24fd00000000,
103'h34c5fb2a5c7ca2fb5200000000,
103'h0ce6917a4f0ae55212f77abd2f,
103'h0b714ff902d0e07c6e00000171,
103'h1c48ab3bceb771f6bc00000000,
103'h2ec044a39928c1efbe00000000,
103'h1cb48106b6716d2b8c00000000,
103'h18b3a2bbe531b1cf2600000000,
103'h1683a4ed82e632d5dc00000000,
103'h240b1915da99d591c000000000,
103'h0abb4f2df21d7a7f422ed3cb7c,
103'h26dcf271972893951e00000000,
103'h2730478460e3e2c31000000000,
103'h2b69cf6d06c0d534a600000000,
103'h083d2ce76cf11cb90666182f35,
103'h182e04e1175aec260c00000000,
103'h3e47706fde98190d7800000000,
103'h0444bec1b6c61dee9000000001,
103'h1002e248340d8e5e6efaa9f4e3,
103'h08b22287b9524d2026f037d3cf,
103'h18bc4eed48552f685a00000000,
103'h095e9460530751f0142ce2c823,
103'h2ec6f7c1eac3a0dd5c00000000,
103'h083ce981f222353dae0f6e5e2e,
103'h1c05286220e92cff9a00000000,
103'h3b2296aaaa2616818c00000000,
103'h284756e3472b3ee3ae00000000,
103'h022fb7f9414dd58e58bfca0000,
103'h113a4e4cea952c719e5290eda6,
103'h3e2e11a02cc4e46ae000000000,
103'h1647eb74fcff32b7ca00000000,
103'h348d042d7a2d4457f600000000,
103'h141ff27451752fccf400000000,
103'h1f480d2cc60233fa6e00000000,
103'h16350c501b22266ec000000000,
103'h0b213e2b3b6a339b861213e2b3,
103'h393ab45e509f3feba100000000,
103'h38c95a5e5ac07e16da00000000,
103'h3e5a3458d2fb32752a00000000,
103'h210d34c20cc48cd38400000000,
103'h3a2a68c6cb1ec12c5900000000,
103'h26e6dcb72b2bf5ee6400000000,
103'h2b63cebe66565eb52e00000000,
103'h02dbf33acd3d3b6c5a33acc000,
103'h2618a48ab6a10a2ac000000000,
103'h17741706fb7cfd658c00000000,
103'h30fb7f71a095a1f04200000000,
103'h30d946917609b8f73c00000000,
103'h3cf4491da7053868df00000000,
103'h3eb055d496de7efa5400000000,
103'h3ce95ff112d2c817fc00000000,
103'h1ab80bfdd2831dec92002e02ff,
103'h2e907101cf6c7ddda600000000,
103'h2b6e0e6ea92489db7800000000,
103'h3e2a2ad5d6b4fadd4600000000,
103'h24b90f550323094bee00000000,
103'h1ccb11c0c04d3421c400000000,
103'h2349920a24064376c600000000,
103'h10ec9c2f00d15537860da37bbd,
103'h1544a131221ae741aa00000000,
103'h1cbfaf7f32078370aa00000000,
103'h2287f1ef064c24a1cc00000000,
103'h0e5677d5a20bd420fe012a0051,
103'h38f652f3c693c6100600000000,
103'h06b1155394ea3de5a800000001,
103'h04735b240ce090d96e00000001,
103'h0a81c5965291a62d0220716594,
103'h349c0429990501511000000000,
103'h224a08cce286c6e76200000000,
103'h26e24b55d622cb10fa00000000,
103'h375b1eb83b6cd3ddde00000000,
103'h19659847a04f1f33b400000000,
103'h1575132816aa3debee00000000,
103'h320b54efee0fd6338f00000000,
103'h26c461c8c284e95ba400000000,
103'h16ea427f74903e4b9400000000,
103'h255f4269dc54a0145600000000,
103'h0b7e8040333ee293cc02fd0080,
103'h1ead944a169e24fda800000000,
103'h346191afa11ca53dda00000000,
103'h00a5cd60beca3987f0b8037457,
103'h293ea926352bcb379200000000,
103'h0216677f74d198985033bfba00,
103'h348c4ad65e1041be8400000000,
103'h061ed36b2126a93dfa00000001,
103'h167b9587d4b2f4145800000000,
103'h1c0422dc1ad1c77f7800000000,
103'h175e48c8b34d5d074e00000000,
103'h2ec8b073ce517fe36800000000,
103'h2759c15ce4afc8ac1a00000000,
103'h349dc65a5278791fe800000000,
103'h1eb392d738d23a7ccc00000000,
103'h3916bc5b6e7000d71f00000000,
103'h22cb65c30d2393ae5800000000,
103'h2e2fd7d6c53a5009c600000000,
103'h0e0cc30a6705b5ccd202408421,
103'h26bbe8bad6358da39600000000,
103'h2cdb0f42654250adfe00000000,
103'h3f1dc9784afe3968d500000000,
103'h149ad3b7f6d948ab3800000000,
103'h131d93c474f712238200000000,
103'h26d5e1748891e5db7800000000,
103'h1ed07fd29caf799fec00000000,
103'h20c9579982855b147400000000,
103'h189b780ba255dae71000000000,
103'h0464aaa1431f32809400000000,
103'h3abfc3125cbaaa8c3700000000,
103'h0aca5523601f552d7800000006,
103'h1e5a4248dadf183fd400000000,
103'h15400a5566a96d633600000000,
103'h0e4504e28403afac1000825000,
103'h2304a9fbda43ba017600000000,
103'h18e3a442a888bee3fc00000000,
103'h2aa1b6c94a8d68dfd600000000,
103'h210936b325710d227e00000000,
103'h1d7466490e12c3ebc800000000,
103'h32234fe06e1bfa9eed00000000,
103'h315af85bcc9060e7fa00000000,
103'h3a2009b6feb3b0c86a00000000,
103'h27562834b10ea9243600000000,
103'h229f0a9e2a2eb2db3400000000,
103'h0c03e7a69084db0fe443ffd7fa,
103'h02f92596f223e5ae0e4965bc80,
103'h36a2144fbf27cd54a000000000,
103'h1c59ac2cc020f2eb9200000000,
103'h2b3ff6e4f8c3073b5200000000,
103'h0aab1cad141cb36812002ac72b,
103'h1e3a28233e5caa4d0a00000000,
103'h30f100ee0a07c6fa1e00000000,
103'h02c8cca46941ef1d5e291a0000,
103'h0f639f961932f00b6891480104,
103'h2c1b25efdafbbcafd000000000,
103'h0a2f5696a95f5c45e80000017a,
103'h334b4e37967a8235c300000000,
103'h02a934f5e0a9d8cc6cbc000000,
103'h2b3a0bbf94f527040200000000,
103'h2ec69f39169e5bf9e200000000,
103'h1ab28ef882d867b9760000000b,
103'h1d1900edb09f06f28e00000000,
103'h3f294baf4b5195eb1000000000,
103'h372ebd74e76a96d8c000000000,
103'h04d28b346493e2880a00000000,
103'h144ec0ad5ac29ffcf000000000,
103'h1469fd18de952b315400000000,
103'h1ed6cf6f72e3ebdeb000000000,
103'h0eae389ec64de8f78e06144b43,
103'h221984562524b8670200000000,
103'h1247700a72d2f105c800000000,
103'h230a86f016ec755bee00000000,
103'h24b189b46833e5666000000000,
103'h2ca675704a3e6c567600000000,
103'h1ac019932eeff60ae00000600c,
103'h3cacaebbdc966b7b2a00000000,
103'h3285b9407756850e5b00000000,
103'h1292a92b730333ca3600000000,
103'h3ede056ce688ed0aad00000000,
103'h181957b9391b96362000000000,
103'h0eeb1580b6f99ba3067488c003,
103'h3a1358568e12f35c3f00000000,
103'h1a3ecef69cfe08dcf600000003,
103'h20f332a1581161338400000000,
103'h20c32c823350302a2200000000,
103'h168cc206154362cb7a00000000,
103'h1b694ae634068f4dacfffffed2,
103'h3d43dca34a935153c000000000,
103'h362fcf93e4fc9c39f400000000,
103'h256bf2aea24078dd3e00000000,
103'h24eb7894d97048712400000000,
103'h1a718dc8bcdc3b1fc60718dc8b,
103'h188af45062c7b3b49e00000000,
103'h3ca0f711fd39417d5d00000000,
103'h02f772b0d4c435cdbe00000000,
103'h22be36c0d3652cdfba00000000,
103'h3e6135f0945c9f908f00000000,
103'h3ccbe8d4f61ad6516000000000,
103'h366fdd36b57c0c41f600000000,
103'h04d807663047f516ec00000000,
103'h26a55e7566b7d24da200000000,
103'h1ccf55152c8fd9b3d200000000,
103'h09142206533538293a108d17b4,
103'h2ad4fb396f048d3e6600000000,
103'h3eddc9837718af44b800000000,
103'h389e6a1b22edaa7e2700000000,
103'h1eeee466a0cb74019c00000000,
103'h177496db5869de1cbe00000000,
103'h3cfed68e7658c2835e00000000,
103'h18a1c5864ccd595eb600000000,
103'h19325efc48cc2fed2c00000000,
103'h368e6c73e06df5737800000000,
103'h2e54580838a0546fc000000000,
103'h1b73061ff12ec0e3a2ffffdcc1,
103'h155f0d965e8318ebda00000000,
103'h141744f9f8f61f0bca00000000,
103'h363d71d10c552ca22800000000,
103'h1303f317e36c719c2200000000,
103'h1cf9354258a9e36d2e00000000,
103'h06719058aaadd6851000000001,
103'h28e00a7ac8a70bc76a00000000,
103'h16a3b13f0e189c201400000000,
103'h28d3c99f76f8a69adc00000000,
103'h12adc56d0c9c57d9ea00000000,
103'h263597bfb47021796000000000,
103'h046475d9c71de6e66e00000000,
103'h2eabf013ee537ea62200000000,
103'h10ec10e8f2b7f47fea1a0e3484,
103'h3ec88997e163e493d800000000,
103'h201523c0314ff57cca00000000,
103'h0a7fa4ceee187f14aa000001fe,
103'h233da483d12da2d4dc00000000,
103'h2cb398b89aad47a3ca00000000,
103'h188d71813eeaec279a00000000,
103'h34b73fc6aa9e84e03600000000,
103'h3ef98d20c32bf6617400000000,
103'h1a697d4fb6e336281e0000697d,
103'h1086b52276dcc348e2d4f8ecca,
103'h048ed91cd04640989800000000,
103'h233581f760ccf5bb0e00000000,
103'h05082133645bced7de00000001,
103'h1ebdf697869150cf3e00000000,
103'h2d508f448c997202a200000000,
103'h0d29688a2b57689a2abfb44d15,
103'h0acf378ad6a7f7deb60000000c,
103'h2ed0d56362d16068e000000000,
103'h1963c40b2ea097f3b600000000,
103'h0e9024b59d716d571a08120a8c,
103'h2f13edfa34d531624800000000,
103'h253faf1d83655617e400000000,
103'h3f3cd0a9b17944121800000000,
103'h06da8a2994b8f32f9a00000000,
103'h2ae9b10094f5c3d94a00000000,
103'h02ce0939dad04e02de4e768000,
103'h1d17b78b06b9ff037200000000,
103'h26daa9ee4888083d4e00000000,
103'h07568f81269fbfc85400000000,
103'h38c838ed4c7a69b69c00000000,
103'h060a305c52d0f937c200000001,
103'h1b0626cecc99322510ff831367,
103'h388a257e92a362816300000000,
103'h3aade3f6aea989502f00000000,
103'h0b4c0c256733aecec253030959,
103'h2ebb2d8be0e192c57000000000,
103'h1cc381176d2d9eead600000000,
103'h1f6f37245ae8cc76b600000000,
103'h0ec4768176ac4d8e2242224011,
103'h254d64ad561b84b27c00000000,
103'h1cb7e59ea4dffb33f400000000,
103'h3f50057acb2d5fe14b00000000,
103'h3cd0f1cda6e5457fef00000000,
103'h30fe2baea4354afab800000000,
103'h3a46ea4220063cc85f00000000,
103'h286fa409910468770400000000,
103'h22c5bdb24a4b52b92400000000,
103'h01011cdaf4baf6c2b6de09ced5,
103'h0571c6fe5680b4750000000001,
103'h2ae8adea1681d14ff400000000,
103'h2163fd4cdcf3984e4a00000000,
103'h212a9f68c6dc46386200000000,
103'h16ac3847674043853e00000000,
103'h20ae859b076ae2ee0400000000,
103'h0232a43e9d171b356ae9c00000,
103'h00aa5b307ec5a0d070b7fe0077,
103'h04fe585ac0f8450f0e00000000,
103'h2e92990a42a2a03f8c00000000,
103'h2091bca7c6a0f89a4c00000000,
103'h2ea7fb7ab63391a48e00000000,
103'h3a83db1e16c54e4c5600000000,
103'h0757ffd0856d49c70c00000001,
103'h16cec4c27ef124e52200000000,
103'h2ce6824ec54924b5a600000000,
103'h3831d17f9b17e9782400000000,
103'h1a426efcc6fe6bc6e800000213,
103'h00c05640ff303d4684f849c3c1,
103'h242f626a5872ac434a00000000,
103'h0ce79349593302844afbc9e6ad,
103'h10b7ada07c6264eea22aa458ed,
103'h1c8633be8b49f837fc00000000,
103'h2684f7231a01a5d87800000000,
103'h08f666caf687d9970238dfaefa,
103'h049ad8f71d0cd0ba1e00000000,
103'h3ea1b011e60337851500000000,
103'h00f27f64aa9e107c32c847f06e,
103'h1e44f48fe93fc08e1800000000,
103'h351f43522a323ff2c200000000,
103'h260662ce89773482ac00000000,
103'h3ef0b9cffc9677d4d700000000,
103'h0079214da29cdaa35e8afdf880,
103'h2c414959608d94735c00000000,
103'h033bb157e206b5c0fe80000000,
103'h22ad4dd90f47ff1a6000000000,
103'h3eb5622f1283b0724300000000,
103'h3d5a51287430fe4b5000000000,
103'h1c8cd49532e6607a6200000000,
103'h1ec60dc2ee40b1a2d600000000,
103'h3147460b0ccd86380800000000,
103'h124c2ec56a9393faf800000000,
103'h2a8215cb1adada060400000000,
103'h329e5d4b2e2708cb6f00000000,
103'h2afb566e18a91e968a00000000,
103'h2e25d5c90b477be1b800000000,
103'h1ee3e91ef742d24fd000000000,
103'h287cd67ae468a818da00000000,
103'h203ccca2424c9137d000000000,
103'h30a5e1602ac967b2b600000000,
103'h0a5671ffca063454f800000002,
103'h1c49d4ef3aac15b52400000000,
103'h12a5dff7860287b4ee00000000,
103'h0b4e7c37a34c5ca42a00000539,
103'h2ec0802a74f23c9bb000000000,
103'h1e38b8723f40b8d35200000000,
103'h095d066f2f0138fdc62e1f4974,
103'h3883dc210c39f1700400000000,
103'h0af70e771496f7df320000003d,
103'h115c7d68cc1ad4003ea0d4b447,
103'h1502a52dd611e2775200000000,
103'h08aa05f0a66e5fe01e622d085c,
103'h068b58237a71050df400000000,
103'h1a03a235821b0afe9a00000e88,
103'h3896c047caa663221700000000,
103'h2f3bc0d164aa05579800000000,
103'h084f213b1c40c59f6207f2523f,
103'h1ed386b2ca7c8670c600000000,
103'h3972f72914cba7abe500000000,
103'h1ab8cac1729f2e5eae000000b8,
103'h22a8a3b16a122587c200000000,
103'h06d94240c6caf0493600000000,
103'h34866740e87393faa000000000,
103'h38ff33ecee4cd63b6600000000,
103'h2e172ef7a2d33d7c4e00000000,
103'h0e414f8a1ad271693c2020840c,
103'h36366065c8e9a060e000000000,
103'h049f053c182aefeafa00000000,
103'h0354804dcf615050c4a9009b9c,
103'h22dd38dbd300558cdc00000000,
103'h1c3862d31554d5daaa00000000,
103'h207d2d2b36320eb67c00000000,
103'h3cece76e556a71899300000000,
103'h26bdf20234e79eb4c800000000,
103'h248f5222f2d486231c00000000,
103'h36b5881e589278255200000000,
103'h3e0dccd03d21ca484400000000,
103'h1cd0830bb2d752669c00000000,
103'h2f7ad7fbf2e51f36da00000000,
103'h32f9b30f4eb5a2428d00000000,
103'h0f0b0647fc307a3e7e0001033e,
103'h293e23c8ee2a2d4dcc00000000,
103'h364893b07c353395c800000000,
103'h353822cee673575eb600000000,
103'h02dd542fdcbbeb0f34b8000000,
103'h0ab2ffcf50f40dde1a0002cbff,
103'h02b2d8bc92d1620df648000000,
103'h36e7e53f9e8461dd4600000000,
103'h1090492161373a99daac8743c3,
103'h06f49812571f1fd97800000001,
103'h0d4cf4e166af68fad8f7fe7dff,
103'h2776b3be6ca4010d2e00000000,
103'h1e24d478b8f0f5ee9400000000,
103'h370a2fcce167a9ad0000000000,
103'h240eaafa7e8c7e25b800000000,
103'h38c28f22f696adf29800000000,
103'h381a74589aa558ed1900000000,
103'h33634f7cd567e8100f00000000,
103'h0a13d44e0c825c68a80000009e,
103'h2250d744fee5abe57c00000000,
103'h3124882e8af980338a00000000,
103'h1a9d92052c4a57788804ec9029,
103'h177e83ebde6edfa71200000000,
103'h20e1d23b390c71ac4000000000,
103'h2a2acc700e8af5981e00000000,
103'h3d6d46d8716cc7d35600000000,
103'h3cfa18b95a9794436400000000,
103'h1af5ca415604db1bd4001eb948,
103'h30fded7594fef3d52e00000000,
103'h16910641eef4be168600000000,
103'h2a90e6e1a0f2ab8c1a00000000,
103'h1b285bc4b683b1ce08f942de25,
103'h20c4abc3a01498afa800000000,
103'h3a5fef97ba3cf4745f00000000,
103'h02eff1825b01a0380077f8c12d,
103'h2c729ef914618fcfba00000000,
103'h0b78fe3dd95181521600178fe3,
103'h0a93f63244c4204b2a0000024f,
103'h06ebe29b0e3d1e890200000000,
103'h1d456f3bdad114bb4600000000,
103'h07008bac60bcf7565600000000,
103'h0b0d296efd0266923000000086,
103'h10dde77cc302f23e90ed7a9f19,
103'h26ebc4138d101bad8c00000000,
103'h16cab5659eee032a4e00000000,
103'h26669e0e04d9c73ddc00000000,
103'h3304ed489ca47ca37b00000000,
103'h02a62ec1c20b1ab17e80000000,
103'h1f578be8761007fa1a00000000,
103'h18f6ec3978b636bbde00000000,
103'h177013c8570dc2a45400000000,
103'h328db7faaf04aeddcd00000000,
103'h10b676de8574c2a622a0da1c31,
103'h24ef3dbc77027aa0d000000000,
103'h30de3b5646b8f17f5400000000,
103'h12dafb946aa82f3bcc00000000,
103'h22dc6ab05a866a921200000000,
103'h36529c726d6166267e00000000,
103'h02cb48d54e3dd0d6d846aa7000,
103'h16fce6b786906d494600000000,
103'h14d6b3d5885bb61e9400000000,
103'h2c36eb859e589cd61a00000000,
103'h32f8895c332f50aba500000000,
103'h08f7f809a0663c314248e21c71,
103'h2287d400535ec58d7600000000,
103'h067366159b56bd971600000001,
103'h0ab79500fede919768000005bc,
103'h002b14980551f7ad04be862284,
103'h1604d0604f098cae0200000000,
103'h3e3d51b60e34a1460700000000,
103'h02cc90a2e53971a656428b9000,
103'h053a61272476c35c6400000001,
103'h0cfa2958674353ff4afdbdffb7,
103'h22c37e37ad7db5266e00000000,
103'h06c1745cf877de7ed400000000,
103'h10f8dc289a3b5cb6805ebfb90d,
103'h3ea70750a0fcd1137800000000,
103'h14988677f2f5ad3c1200000000,
103'h1407bac5b09cb48cb400000000,
103'h0eeecd9245353b04a612048002,
103'h21113d155a3cf5ca5600000000,
103'h15307dabe92bc35c9c00000000,
103'h3a456b7e893d0071f700000000,
103'h12f70ddddf6d7e1dde00000000,
103'h2eddeb41d8b2e99c6600000000,
103'h2401be702aa9f77a4400000000,
103'h025154fb1887e2bc1e3ec60000,
103'h28ddebf7fc89a12c4800000000,
103'h2ed80112bedaf6276200000000,
103'h0c84ffc9e8b8e21f5e5e7fefff,
103'h14dbf5fb5690e3321e00000000,
103'h36bacee8e315e2fc0600000000,
103'h16234902b6f1d8f75c00000000,
103'h3566b943eeaca7e03e00000000,
103'h3b630ba484cff0e2f400000000,
103'h16f041373836aa26e200000000,
103'h149359c5f299b5cb6600000000,
103'h09284b4c0889f7029ed0de274b,
103'h2d69e4b25c1d50c89000000000,
103'h127b6efba4459c149800000000,
103'h32c3a36bd0af80c6f500000000,
103'h02a58da7652aefc29ada764000,
103'h1d116ee596ee932e6a00000000,
103'h109aa0ec589420d5ce03400b45,
103'h2a696f07b4a58fbb6400000000,
103'h16e7bdea074030a7be00000000,
103'h2490fc8ef0a99faf7200000000,
103'h0a28ce6246915d997800000001,
103'h0954c10b6d225a286a3b4d9183,
103'h3b26436ff64b288ab000000000,
103'h3537f67c3e9fe9961c00000000,
103'h1ef34937f8c62d061200000000,
103'h0e3ff98d2cfe2382501f10c000,
103'h2caf040acaf16cba4a00000000,
103'h3f6937131a3166477700000000,
103'h10c353b186e06a5242f174afa2,
103'h1ae39d560549a1655c0001c73a,
103'h10020a7cd50cf516e27a8ab2f9,
103'h1211e45deef0926ce600000000,
103'h2f53248680f29ce9bc00000000,
103'h1074cf0152048147aa3826dcd4,
103'h38e01ae18257a5ce2a00000000,
103'h34585bd892cc74cf7e00000000,
103'h1ec12f3c8aac8fb10000000000,
103'h0a1c9f8a3e04eb8992000727e2,
103'h097c911f9ec61ac61edd45ecc0,
103'h0934288328e2ba505ceb4969ba,
103'h1ab834b6305f4b6ffa00000002,
103'h38e8d09a389373f32200000000,
103'h161e5807d24ba8a95200000000,
103'h1119fa3b8c3479438a72c07c01,
103'h34f856bfa352d14b5e00000000,
103'h0635feb3b36ccb86ea00000001,
103'h12071a9ae76522468c00000000,
103'h3123df2b6e9b20fa3e00000000,
103'h1b751cff80a23b9526fffff751,
103'h27192c1ef0c61ac09400000000,
103'h252a06c54b3b37c01400000000,
103'h0aa003b2315463df0414007646,
103'h1eb12199557e6aa44e00000000,
103'h33647b15a11e6e567f00000000,
103'h36ddef527ecf8fefd200000000,
103'h04929b4f72340b057200000000,
103'h029bab2b6911fa57f268000000,
103'h172325abaea495a76400000000,
103'h08c90e82704040d2cc44a7285e,
103'h3a3e87490663667e7a00000000,
103'h1ee80b15112c7500ec00000000,
103'h2ca389390a6afc49f200000000,
103'h27039d046a53075f0200000000,
103'h12a3f1a296f690980e00000000,
103'h06a7acbf3cfa2d9c7800000001,
103'h08d7dcdcd09e1f3f0e24e1f1ef,
103'h177309445645cbfe4a00000000,
103'h0e613d0ade1da8db1a0094050d,
103'h1d4601697690b21f7000000000,
103'h2824f36484f1ef2a5000000000,
103'h02a2049ea337f093c688127a88,
103'h3564e1d70a5ce3f84a00000000,
103'h044567ea8cfee896ec00000001,
103'h0ab6a01d8063ca6df60000000b,
103'h1419c77ac4a932588400000000,
103'h02b4df6bce5fd2760469bed79c,
103'h38acdb55257999f0ca00000000,
103'h3ca3bfd5662e795c9800000000,
103'h02fe6ec39edb54b1bcc0000000,
103'h0d02500a5c7f148722bfaa47bf,
103'h256603c71f7d834ac200000000,
103'h23435174ab7fd3551e00000000,
103'h044f187ecee5d71c3c00000001,
103'h0636343ab1292890e600000001,
103'h249c647db678410fb400000000,
103'h2080180b7cae754a6600000000,
103'h06e39eee634ad9c81c00000001,
103'h3c2cfced82caf1d39900000000,
103'h229f837d8aae90c1fa00000000,
103'h3e8a4b1d46db8daf7e00000000,
103'h17238807697b112d0800000000,
103'h13079eb9a7055c4a4e00000000,
103'h10b6a73f7d28e451b6c6e176e3,
103'h181440874f30830b5c00000000,
103'h264d677e9ee72a4ad800000000,
103'h1c019fa2f6fb6ad22800000000,
103'h38bb34119c48d250c600000000,
103'h109dacd1f94a71f3bea99d6f1d,
103'h38b0a89db005a6055a00000000,
103'h00aaceb442a352d754a710c5cb,
103'h3ea05f9cfa53fb750500000000,
103'h18dec2d67afeca294600000000,
103'h2c679803b89f29c64200000000,
103'h32f61336527dec9cbd00000000,
103'h3827e1403ee584a07700000000,
103'h3aadaabf30db97d6c800000000,
103'h39323e676a0379170700000000,
103'h2e55fbd5e4b123d63800000000,
103'h36f7a5e11ce3623da200000000,
103'h3c7ed48cca395e138600000000,
103'h34e19b0f413103f4a400000000,
103'h1747daa8beafd8816e00000000,
103'h1e5f3e1872917390b000000000,
103'h035a03c5cad94e396e72800000,
103'h308e2786a8388c51e000000000,
103'h20f34f3c2a929017aa00000000,
103'h0e084f731a20b79e5200038909,
103'h30aec33abc1406da7c00000000,
103'h1a2e853bcb1c564d9800017429,
103'h2ee6d38ebacb19885400000000,
103'h2b31b1f956f99ec41e00000000,
103'h029d480244e07252da80244000,
103'h161ce4e5af12244c3000000000,
103'h36b8d816b2af6c4e7400000000,
103'h101fe4d008cc513422a9c9cdf3,
103'h0080904d7e85294ad482dccc29,
103'h34c1ae1dcea50e1ade00000000,
103'h1614f03a4e259e685c00000000,
103'h2c179ea542e74c862c00000000,
103'h0ae69e445afc3cc07a00000003,
103'h273ac72e4713db65be00000000,
103'h1333fe3310fa79aa1800000000,
103'h0e52d3a0373540d85e0820400b,
103'h0d58f5938b693f0b6ebcffcdf7,
103'h255b544758bc12aba400000000,
103'h03718e60e415083f2e39000000,
103'h3082422488705c868600000000,
103'h14c836c08ae1eae76a00000000,
103'h05776a67fa642d0bf200000001,
103'h0ae2b0bb0e2c63cc7c00000001,
103'h3662ff4d52a3ce347600000000,
103'h2953aa661e867eef8600000000,
103'h2726406654e97e3cd800000000,
103'h1c5d03727c3d28a2f600000000,
103'h22c02a4b226369094a00000000,
103'h3cc71f5840c06c7bc800000000,
103'h32549354e28096c6eb00000000,
103'h3ecb858e5e47b61f2b00000000,
103'h077fa06ad29c49740e00000000,
103'h309724509067cf026c00000000,
103'h1d6f14b216e76f6d3e00000000,
103'h2ac79bda867e93bdce00000000,
103'h1667d92222eda86fe400000000,
103'h16a45fddccb5444a6c00000000,
103'h2548b59be41d1d6c8e00000000,
103'h0ad47ac73ac17d4a5c0001a8f5,
103'h36ded3b05f0a32e64000000000,
103'h04d6d50968deadad7a00000001,
103'h20841aacdebd815dd800000000,
103'h214e7dbce49456674200000000,
103'h1ada5e17441871142000006d2f,
103'h35707157e666eed10400000000,
103'h36e5324601414ce84a00000000,
103'h16177491f4b1be403000000000,
103'h1cde0d452a96f0863000000000,
103'h26bd170c82ae65182600000000,
103'h17030fa4de8c725d5000000000,
103'h068a552584498969d200000000,
103'h2cc358e65a4c990eb000000000,
103'h3e934d2d60d6ee343400000000,
103'h1111a68c8e9a471a8e3bafb900,
103'h031c72490d2d9447f086000000,
103'h3670c76f5d3f3ad47e00000000,
103'h0611b5a45f5bad1d8a00000001,
103'h3689920d96cc748ce600000000,
103'h349bb5915cde2a314600000000,
103'h3edb6d5d1367bc3edc00000000,
103'h255a5ffd470371d03800000000,
103'h2b34ffbb04dedf2d4a00000000,
103'h06dc1405a9393f2a9000000001,
103'h3f615281956e3ee59400000000,
103'h084e4d3c5a4a52eb3c020febb3,
103'h193eb9c75aaba56cd000000000,
103'h2c0e057fa2f9f2a92c00000000,
103'h2b1690627d38ac708600000000,
103'h3a8d5a2ae846b1f02900000000,
103'h264e76de925d4252a400000000,
103'h2cbb38ff0eea9c7d8e00000000,
103'h1621edc8b439135c2000000000,
103'h3ac14f02e2f44c5b2e00000000,
103'h08a7622d39163a23e4d8ac076e,
103'h2aeab7aa32d78926c600000000,
103'h1918a9a4bd7eeb53fe00000000,
103'h3d7faefb6669a2fe3000000000,
103'h02db00ad3e824ca2eca7c00000,
103'h014c8c82fc01fb9e52a74410a7,
103'h3295a17f7edcfc4b9300000000,
103'h1f5da1d0012988ce8e00000000,
103'h328f451eb2bf2a4e0d00000000,
103'h04433510501ccc1e0c00000000,
103'h12f920a042ac113cbe00000000,
103'h1e8c087bc6ef464d1000000000,
103'h2c487925d8e866ed5200000000,
103'h2ac4141df9746f691a00000000,
103'h3b5c7b3424bce88ef200000000,
103'h0ea0f3870e80fcacea40784205,
103'h28d4b2270add77e10e00000000,
103'h1af0d7b4597e6b681e0000f0d7,
103'h06816caac1531d8f2800000001,
103'h14ceea301b43f5438000000000,
103'h329d646260c561ee4100000000,
103'h1b495675b6944c1e5afffd2559,
103'h1a73b3f12931b080bc00000000,
103'h1af12efbc57b06f6720000003c,
103'h36b29f49deeebae79a00000000,
103'h333971863adfe9e35f00000000,
103'h25548fe0f092892d3e00000000,
103'h3ea15ebc62cbfab37800000000,
103'h1f69348e47208a946800000000,
103'h1c1fc547c4c1e950ca00000000,
103'h14b63fe4a32b1ddf1000000000,
103'h3cdf43aebe4ae326d400000000,
103'h06d4422c5301230b7800000001,
103'h16e9cb3e4ee066ba3600000000,
103'h2ac13da114b4a8e68a00000000,
103'h22c3cde2ea9e7424d800000000,
103'h1b11414b975fb1c5eeffffff11,
103'h245fd7bfb8237fa8d800000000,
103'h3c8ed4ee1234c0f46e00000000,
103'h2a727b02f69498b42800000000,
103'h04f4953cb4236da23a00000000,
103'h32d6613c5e95e8a53300000000,
103'h1adbace4e28a7de1e600000dba,
103'h1715b981d660df1e4400000000,
103'h08e45ed2f13c8c0328ec6968ec,
103'h2ed671c647524584fe00000000,
103'h325e6d5ece36a457ef00000000,
103'h1a70e6d93d0d161e3600000007,
103'h18e43f71f06b837d0400000000,
103'h0894240dcadc6a564224272dc4,
103'h3e964e2ea4c0a9c83200000000,
103'h02cf1ca76c54cdd5fc80000000,
103'h0515013e6aeb1c04a000000001,
103'h36c669526cba38ac0c00000000,
103'h35543bbcb2cf39ea7600000000,
103'h14a2b7ef2895a33ce400000000,
103'h224601f79ce9def99600000000,
103'h18d46804b28c96e8be00000000,
103'h3d1d06bdd4d298e05c00000000,
103'h1234df616ca700e50e00000000,
103'h12e25b41eac407a2e200000000,
103'h2e79b61bfcf8e7044e00000000,
103'h3c9da7decedb42463900000000,
103'h1e943281fd54f8623600000000,
103'h2c31be0a38f2a0410400000000,
103'h269351355686d2c30200000000,
103'h1cedcb64c4b890cd3a00000000,
103'h212387da6b4be2029200000000,
103'h22ae3cb24739ad675600000000,
103'h1e2b91cb275d3541c000000000,
103'h312fb9a70b0b71f40600000000,
103'h06ec7250283703bf2c00000000,
103'h06f50cfbd866bd663600000000,
103'h0d37550ede532fb65ebbbfdf6f,
103'h38d6d263a4483cb23600000000,
103'h3081c1ac707f91c11400000000,
103'h0e63b4b468566424b821121214,
103'h06ac652298d825d12800000001,
103'h1b484547293bda8592ffd21151,
103'h152c621deee83fa82a00000000,
103'h3c9010b5c83084ef5200000000,
103'h0e4a23725c5ce70d4024118020,
103'h3adc5c001aecf7c30a00000000,
103'h0caa6f1368371b35665fbf9bb7,
103'h0e60c1cee21377358000208240,
103'h19479979b0bde648ea00000000,
103'h3e8b5831be1ea817cd00000000,
103'h00bc0eacd66641917c91281f29,
103'h2a23e05d54f199c33a00000000,
103'h369f294354ada8701000000000,
103'h34d858723ed188cd6600000000,
103'h2f302fb8f670b210ba00000000,
103'h00ee48912b490a82fa1ba98a12,
103'h269dfb2c99793a3bf000000000,
103'h20fb5638196782cd1a00000000,
103'h1a2a3a10fe057df9b20000000a,
103'h0ac9cffaa100d431cc01939ff5,
103'h24b270673a2b0e42ca00000000,
103'h19144b0fc6f4de3d6a00000000,
103'h24dda8856aa74ea4a600000000,
103'h2eac83f4c2bb99b46c00000000,
103'h1a7c3395e6994239d60007c339,
103'h0176f179d745c62e9a5e5bd438,
103'h2d668d9b30c1f9c48000000000,
103'h02fd78613038eb3e56e184c000,
103'h1d4ffcdb9c9f78d98600000000,
103'h1e3bc38fde9cf13ab600000000,
103'h356d5072bcecee165200000000,
103'h3d60d71a1b28b1a63200000000,
103'h328d48ffce960218ef00000000,
103'h065933bf0af6d9330800000001,
103'h38c20fb8fe842232d600000000,
103'h2717d9c944dd55f1e200000000,
103'h2e96557fbc9f65aae000000000,
103'h04aad34f22b73f742400000001,
103'h26b62a51914d94f3e000000000,
103'h0645a386d4f868430200000001,
103'h2ab272adfcae92949200000000,
103'h0abea78002f4361b6600000bea,
103'h0c821bc62ea6a8c962535de7b7,
103'h1e932500396550496600000000,
103'h069c967d46e76c0f9400000001,
103'h28549a8ee47a910fcc00000000,
103'h0e00d4bbea17278d1200024481,
103'h2353b7b2556bc21bf800000000,
103'h300beaf2226c96d7e200000000,
103'h02ab8a4186c04e8a3618000000,
103'h3ac5baa0b6cc397c5a00000000,
103'h1ef7128cf977c3bde000000000,
103'h14942c95353d7e5e9600000000,
103'h2e9ddd75523490eb8e00000000,
103'h0e67dcdfa6c8bd80c2204e4041,
103'h24fe15c656669af61400000000,
103'h340c126ae4ce77d5bc00000000,
103'h37578d6e0acc8d9c1200000000,
103'h0cd7995cbed8a006f66fdcaf7f,
103'h082062cc34302d75000827dc9a,
103'h1acfc731c007c6d1be00000000,
103'h104da36d0928299df492bce78a,
103'h12980d4462f7f0cfb400000000,
103'h10bb1722b545943cbebac172fb,
103'h050e4e7606dda1812000000001,
103'h3a694c9b1698b8a3d400000000,
103'h38ec745e1ca70719da00000000,
103'h19678cf0d71053b4f200000000,
103'h2f2839c04efcc8130e00000000,
103'h08c68810e7645503e4d16e8981,
103'h3afd8f05548c8ec43300000000,
103'h08db9d139e5316d5184445e343,
103'h2cc9fed6d950a5da6e00000000,
103'h1eb528ad232c42ee0c00000000,
103'h3804a7874ef641c4e500000000,
103'h26e0b525aeab6a720600000000,
103'h330fd99926b011f95700000000,
103'h168fa3e70c90c71f0400000000,
103'h1f3bb122fea0a0b82a00000000,
103'h34de0023d530449f3600000000,
103'h382bb996b36bf5c23400000000,
103'h22298502e649f5e60800000000,
103'h18b8178e1f75af7cbc00000000,
103'h0ce74ad1809f347fa27fbf7fd1,
103'h1446c2b419574c0dc200000000,
103'h10123058e43e96df42e9ccbcd1,
103'h352793e3ba8559935c00000000,
103'h36b2a6eb4a9789ec4000000000,
103'h38dcee727ebf1dcffa00000000,
103'h145e82077571c4bb4600000000,
103'h171eac7bae4eb32dc400000000,
103'h1064308342ad35353adb7da704,
103'h16413e7718cbe1b0e800000000,
103'h1cdd6a3aea3012342a00000000,
103'h16eb5aba017150ab4400000000,
103'h3e47fe66dd4ebae62e00000000,
103'h2851d748f23a15a02e00000000,
103'h2c2791dbf08214070c00000000,
103'h1b2d5ea31ad3eb4ffeffffffff,
103'h0aa47c1586fb7d2bf000000052,
103'h176a546e2328dbcf0a00000000,
103'h156a4266eccd57e49000000000,
103'h04ec4466c237ac52b200000000,
103'h0e4231b696a1eeb99e0010584b,
103'h20939c325c8e33206000000000,
103'h120de27d2ad064d6f800000000,
103'h325580ac8b6401095500000000,
103'h12d4cb2e9e71e3867e00000000,
103'h0af6046a50c764330a03d811a9,
103'h1ea570c6629c2f61a800000000,
103'h1f2541f96e9233cbf800000000,
103'h28091435cc37a4925a00000000,
103'h105ec9f8aa5ce68bc800f1b671,
103'h087be3ee9365fac1968f0c9782,
103'h22352d4622c4c4ba4000000000,
103'h2c80aa69ab40a8a8d400000000,
103'h0303cc1f8e75d5eef638000000,
103'h02e3d4613af68058a2613a0000,
103'h1729d7647cfa4c783000000000,
103'h0e349f21fede20d96a0a0000b5,
103'h30800f885707f83de600000000,
103'h214155dda43c975fe400000000,
103'h0af91c8b94bca6e83a00000003,
103'h30ab2fb1b4fdfcc5de00000000,
103'h153b63b13ef719517200000000,
103'h10d38feeaea249032618a375c4,
103'h2ea8538c02ddacb46400000000,
103'h2239be1192b13ca31200000000,
103'h08c9255d0359902f16c85ab90a,
103'h2f4fa5f9e4934e40a800000000,
103'h00786f99ec5c739daa6a719bcb,
103'h167ee5ee5aac19978e00000000,
103'h013698e5dd2489317c2d910bac,
103'h2a47dc0c72a36f1fd600000000,
103'h3aec6d73b2da0805b300000000,
103'h36ed72789f21e4122600000000,
103'h0c9a9115180e5185d84f68caec,
103'h016c38e30efbc3fe7633fe70c2,
103'h26e14fd0da9655138e00000000,
103'h3e306ec45a028df69d00000000,
103'h36a171ca00e3ddc77800000000,
103'h0520c65580144c8bd200000001,
103'h229bdedf76b5be55d400000000,
103'h1aad4c7cfad684ab540015a98f,
103'h2cc148111d72638aca00000000,
103'h00b9216cb61fb007c46c68ba3d,
103'h14c5475424e0f818e200000000,
103'h1e872b91649a19859800000000,
103'h251f9479fa5f60d9bc00000000,
103'h062a60ed58e68c6b2200000001,
103'h1e54dd687d0620e51c00000000,
103'h1c6051fc823081d27400000000,
103'h3f05e01622855f3af300000000,
103'h1b0acf097ee5b13774ffffffe1,
103'h0ef64a67fceb914d96710022ca,
103'h00e7e6ab96f6605714ef238155,
103'h360a04c1a4ecaabf1000000000,
103'h0cb18212a6d4916aa67ac9bd53,
103'h233eb09b1cde962c4c00000000,
103'h32b770712890183ef300000000,
103'h1a26909e4acec8da0e0026909e,
103'h26825b8a7e86394b3600000000,
103'h18b2b7e158acc9e98200000000,
103'h26c1aa647f2f25740000000000,
103'h1d60b52696e1dd555800000000,
103'h1ece88c2bca387b9d600000000,
103'h1ec295aa19043ce06c00000000,
103'h37636c7af8d2c5a32800000000,
103'h0c3368bfd6955b4d405bbdffeb,
103'h38e5425a0ef8c7c83900000000,
103'h203aa3ae1b2c30881000000000,
103'h229441e2951172e21e00000000,
103'h1ac0a5ba344c16903800000006,
103'h2a8264df16e05872cc00000000,
103'h093cebcc32a0fe2d02ce0af098,
103'h0223a3415c23630c181a0ae000,
103'h0f1bcd98a6604ed84a00264c01,
103'h11600e802883f219a86e0e3340,
103'h2a84a7da769fbfb24e00000000,
103'h354a3f61c8ffce327600000000,
103'h1d3339f53284760cec00000000,
103'h2a7c8360e6ceb56eb400000000,
103'h2149bee64401ef63e600000000,
103'h0eb6ba1def7e72c4ce1b190267,
103'h0323838810c831ab1283881000,
103'h2b14c2ff1e7eebc90000000000,
103'h38d4b7e4e0a26f511000000000,
103'h0a969c2e8ab732502e00000096,
103'h0ad6f33d028bea3510006b799e,
103'h1cdf7bf68c2286639a00000000,
103'h0b66f07918f979a09e000166f0,
103'h1a90d44cb4d8f5972a00000243,
103'h3671ea707e3fe6104200000000,
103'h14deeac95ad0ba5cf600000000,
103'h3f6e7185d142a4cd7700000000,
103'h02f771e2e5218f96d0b8f17200,
103'h385967d72290011ca100000000,
103'h2efb43dba48772ff8400000000,
103'h3f6dda3d1ee0dad6a700000000,
103'h1e23156c0cdc1eb24c00000000,
103'h22f9e031cd49f8ef6a00000000,
103'h0a60ac142a6d0e5b7600000006,
103'h174eeaf60e66ee8d4200000000,
103'h011e04ae98c79aa16ef2cfa803,
103'h36c93d196f1685977c00000000,
103'h3abe6e73af348a461500000000,
103'h2820ae2964fdc75f8200000000,
103'h24e9dc6c5ebc35d33000000000,
103'h387aa550c6dce3fc9500000000,
103'h3a21f3ccaac6c068f400000000,
103'h2afdcc8ea24165b9ba00000000,
103'h3ed76cb01d6359866600000000,
103'h326d42a4c66126150900000000,
103'h2edffc96073892c52600000000,
103'h141976f038a5d569ec00000000,
103'h1c9457042685d1fff200000000,
103'h0272909e7a9f48f02ccf400000,
103'h30b1f04dd8339ff45200000000,
103'h2229e2c25aa63092ce00000000,
103'h0e47aaa0cb5820e0a620105041,
103'h22eb447f2e8203a30000000000,
103'h302e274dbcc9ae43cc00000000,
103'h16a4aa109eb4f2c2fa00000000,
103'h16c15d664ee31a10b600000000,
103'h2236319ca487c4215600000000,
103'h1d2d0975fc492187a400000000,
103'h14ed8f931f7f53244a00000000,
103'h2b6308733cac5c9a4600000000,
103'h0ebb9b641099ec2d644cc41200,
103'h189bf2763afcf4a0a000000000,
103'h1ec56b1008b89004b000000000,
103'h056e36ce2254827aea00000001,
103'h24c35f268119ed8af400000000,
103'h16b273ac448824591600000000,
103'h009e7cd2aa4b837f9675002920,
103'h354315fdc0fdf72bdc00000000,
103'h0a3c31a3c09c73fe8603c31a3c,
103'h234f3ad4b6df89fc4600000000,
103'h3eea685ec01bbba00700000000,
103'h04d11968626af674bc00000000,
103'h0ab5c19de1555ed37e00000000,
103'h1036ddd1e426783be00832cb02,
103'h0e9784022edc39d9c24a000001,
103'h0d13e5d2801317aba689fbfdd3,
103'h2cfb3e178eaa9badd600000000,
103'h2f37f5301abe81805600000000,
103'h169b248486b9bf97e400000000,
103'h2cda8db2b6f1b4c7fe00000000,
103'h032d0e8c8c8cd94c845a1d1918,
103'h272a2b14386766ff3a00000000,
103'h24e5c91c3a94758bc600000000,
103'h295b26bc20bea09ffe00000000,
103'h24c2392404a469bc3800000000,
103'h2ab624d86cff90785800000000,
103'h2a11778c10c1c99c5c00000000,
103'h23013fcb7d77ee74ca00000000,
103'h3cafa8aae6896600da00000000,
103'h18027b46888aa5cc5600000000,
103'h2254de5a843a4e773c00000000,
103'h3f690b0adf3cc9bdc700000000,
103'h14f526300091a8184a00000000,
103'h120aa755fefab3232800000000,
103'h18aace4854efd9532a00000000,
103'h228543b1e6fa80a92800000000,
103'h0c9c82d93ea54ef17c5ee77cbf,
103'h36456a18e02a92a36200000000,
103'h1ee9047bacc7157ca000000000,
103'h1c7c7831a30c7f958200000000,
103'h3f0a6c90c2f584112f00000000,
103'h213dafe15f71fc42d200000000,
103'h229b85d55d7c68d39400000000,
103'h10c07145fcba18b4f2032c4885,
103'h22f1dc4c1e559e8a4e00000000,
103'h3718cb6371160fd04c00000000,
103'h28b1b6bd9207ec1c6a00000000,
103'h38c70aeb4a20b77fda00000000,
103'h049677cdf2d26e3d6e00000001,
103'h2ebb833aea997928b800000000,
103'h0af69e782e2ff0f6aa000003da,
103'h3939a5d1deeb74319700000000,
103'h309d64ab68e212a9c400000000,
103'h1ad391c2601bb87ba2000034e4,
103'h30a3380210b91d270a00000000,
103'h36a2cf386a8caee96a00000000,
103'h188ddaa05c2fe6eb7a00000000,
103'h255af8b212d2b623e600000000,
103'h0e43cf3f6b6090c44220400221,
103'h0ae5c2f3cebb897654001cb85e,
103'h311465919eff58b5be00000000,
103'h3372ef1ae8e51ba98f00000000,
103'h06a42ec818f9813b2c00000001,
103'h0535ff398b6c70561400000001,
103'h1283592151109f1e2c00000000,
103'h3ed00bbed5469e57b600000000,
103'h1301da05e8c9f7790600000000,
103'h3e2d2988269a0337da00000000,
103'h34c4e9607a9bdd3dc200000000,
103'h3a6d4856f8c906c5ea00000000,
103'h175c45a52e8df0266400000000,
103'h18153a6c68fb387d5c00000000,
103'h0268326b7e577e228a8326b7e0,
103'h275707a8596cb88ef400000000,
103'h040ee3ab1ad4eafa7200000001,
103'h0f54afd4422bf2a2ca00514021,
103'h0295b47ac73ad64de6eb180000,
103'h362e3743d48f86222800000000,
103'h0133729bd9253a9cee2c569c63,
103'h270d98ee4e5371e0c200000000,
103'h0e13b1e38e86e47c9a01503045,
103'h3d54a126b6947d6ae800000000,
103'h0025168c04a82f4e7866a2ed3e,
103'h1b1ac68e42fcd0752effffff1a,
103'h0563e8714221e7013200000001,
103'h3c33eed0dc3cad8f7500000000,
103'h2a98729b60a09600b600000000,
103'h1ca525b45cd484d19400000000,
103'h12aea942866cf76cf400000000,
103'h08da13d1e5121d2152e407785b,
103'h1d422bf0b6c0c663d800000000,
103'h124ada103e9ada35bc00000000,
103'h25280d015cdd06267200000000,
103'h3d72375f6f27e036b200000000,
103'h3ace7eded34fed380f00000000,
103'h2ceb8cc20ec224977c00000000,
103'h1ea374db0890a3764e00000000,
103'h2d38631a767c30385c00000000,
103'h28f53190951fa5136600000000,
103'h3701ed3ec358082ddc00000000,
103'h14d0cd846a4d39be7000000000,
103'h3b305140624f26fd3200000000,
103'h170c0534b71ff4819e00000000,
103'h07075e3c715045c20000000001,
103'h3b5abf72075c4af6b600000000,
103'h18fb5a660d63a9332600000000,
103'h18eb1c5746be68a52c00000000,
103'h0efad2ca1eb9c30b385c61050c,
103'h345acefef6a4df628000000000,
103'h2017162a849fb22c9e00000000,
103'h1837068938fa812b9600000000,
103'h18155f8d181197561a00000000,
103'h38ad7b9c33489ddf5400000000,
103'h0eea770dca5dfd6c6c243a8624,
103'h28c724ac020b79089e00000000,
103'h3c9e5375d0f5f0166b00000000,
103'h2a871995babd14c26c00000000,
103'h08b87d94f75b68383ef18ad664,
103'h3247df00a0e281cdf900000000,
103'h20e2b974ea9aff62ee00000000,
103'h1e7383ff9ce2de639000000000,
103'h16c1634cbcc597d87a00000000,
103'h046aaad21a391bd81600000000,
103'h14f6742570fa7f24d400000000,
103'h0f1d3cdbb66529f6ee02946953,
103'h2626e3f58b5b9e1c6000000000,
103'h3af622e7db78daf81700000000,
103'h28fe7db2409fbeeda000000000,
103'h090157a17a95e1d57aca5b3a00,
103'h1e695b87a2945f87ba00000000,
103'h012cfd8a2c95b72934e15a59b0,
103'h3a697a84caff12b0d800000000,
103'h3645b66d0b2c103b0400000000,
103'h2ab7d42ac6958abfce00000000,
103'h02be51703cdb412cda1703c000,
103'h065a85dee6931557a000000001,
103'h16f5ccfe6b5166c7dc00000000,
103'h30bd2458f0abeca6c200000000,
103'h101a067346a1b9a52cbc26670d,
103'h2c5229ba775eddfe1e00000000,
103'h2e1d62594678e4716400000000,
103'h1c3a01bff2cb0e2bdc00000000,
103'h3b028dcd62e870852200000000,
103'h1f6cd37fff2272451600000000,
103'h3b35f730b92500127900000000,
103'h1e77ff52d691d3927600000000,
103'h348515a0d2c7cac32e00000000,
103'h2d7a9c73f03fca160400000000,
103'h2292958c24c4dfb6d600000000,
103'h10cf8eb6d03f7c2ac648094605,
103'h149e5b73f2d211b6ea00000000,
103'h2d34f2f442a1a06dba00000000,
103'h320b548a963ffbe1ad00000000,
103'h1ea695d7c274eed5ee00000000,
103'h1881534fb68043608600000000,
103'h072e227e9426d9384800000000,
103'h347c921b2ca82c87fe00000000,
103'h3a0afd9972d64f069200000000,
103'h050e57eda952e121c000000001,
103'h0291f5a2625ddebb3262000000,
103'h163c6c8f666c36a8da00000000,
103'h168f10046afe2c4b3e00000000,
103'h08b80280003a98daa4414d2d52,
103'h2533d61d56c9a8df0e00000000,
103'h220d8875de81ab5f0e00000000,
103'h0653717742b5817c6400000001,
103'h169786c3e4c309f24400000000,
103'h251634eb2c167b698600000000,
103'h0b5e8bf182ae022d6c000002bd,
103'h0e288e56e6c437189800030840,
103'h14a81238b122c30a1a00000000,
103'h00eaa00cbe4b5161009af8b6df,
103'h1943a94a54f36399b200000000,
103'h324ab4b554de03a67100000000,
103'h3515f738ee21acf0c400000000,
103'h2603fcc6a16c61a61a00000000,
103'h163d53b5548258df0800000000,
103'h1c6a0e3dba8655a5a800000000,
103'h3774cc6c92c3a95afe00000000,
103'h3ea1378c2e2db798b900000000,
103'h273a0451e4a284054a00000000,
103'h255529f6a243bb917800000000,
103'h1ef6a541087dbfe35c00000000,
103'h295bc9e66ed2e9d9fe00000000,
103'h22eea6248cc98f1b0800000000,
103'h3e240667f52559017600000000,
103'h3e9d223cd713ff260200000000,
103'h0693fdf51638058df600000000,
103'h3d5dc38754d527cace00000000,
103'h3ef118349b6925bfe400000000,
103'h34a9c5e356c6e9473800000000,
103'h037672b814b8017bd272b81400,
103'h267b251ac961c75f2800000000,
103'h1f54ff484cd83a173c00000000,
103'h3097ff35b2535f320400000000,
103'h18a1e86a52a85e7a5000000000,
103'h1463d31ac3405db00400000000,
103'h1a87852a5ce2461a5600087852,
103'h2a837151304619351800000000,
103'h2ed2bcaa0acd9e5f7400000000,
103'h04ca667d37510fb0a600000000,
103'h1e026e006423cc5ab000000000,
103'h131cbb9deaee32d7e600000000,
103'h397d227088f0a0d84d00000000,
103'h2aab27a29b0d5c763600000000,
103'h112a3c85548a7ee6be4fdecf4b,
103'h1ccd1dc2be35a6895800000000,
103'h125e31d80e5fe30eac00000000,
103'h10dfe6c5ac2d00d16a5972fa21,
103'h2a6ef8297e8b32a97a00000000,
103'h16888874116b196f2600000000,
103'h02d7bf47fada1198a48ff40000,
103'h3c86d92a90629a0cb400000000,
103'h2262f3de923a5954ae00000000,
103'h06ca413c0ec1327f4000000000,
103'h3c9ca808b024265dd200000000,
103'h2b49206df8ee6799e200000000,
103'h2b5832dff48b0fa29200000000,
103'h3ea19ea69ed430108a00000000,
103'h20ac3cec8a2c62f07e00000000,
103'h32db019048ce01971f00000000,
103'h3ef82dcde97a3e83a800000000,
103'h3ca069ae1b554013f100000000,
103'h1a1cd59ed94d6de1d80000e6ac,
103'h02c5a48016edd78ff216000000,
103'h323c74f8710aad2ecd00000000,
103'h0b2d83f474d051aee200004b60,
103'h3e73d304660cc6a75300000000,
103'h0b078ff6323a4a9bc61078ff63,
103'h2c892477f0ae1da02e00000000,
103'h3f1566287ab5ad966100000000,
103'h0771f987e73ed20e5000000000,
103'h34db538ea5543836ca00000000,
103'h147ef8312ac631beb000000000,
103'h24d0ba73dea1854d5400000000,
103'h2ed82a4cf3207d7e8000000000,
103'h1e1e6c3456f137f25e00000000,
103'h32b8e65284c9623f5300000000,
103'h3219922f62e7ce73a900000000,
103'h131bc35996a0b4c62e00000000,
103'h243e720248ba46f59000000000,
103'h0c52589d5ad60a4f266b2d6fbf,
103'h3a2fa177bf147c517100000000,
103'h0cf4b8c5cc66d4eeca7b7e77e7,
103'h325a84da069676668b00000000,
103'h227a97e3d28b2f2c5600000000,
103'h2f70b53cc6e5b4065c00000000,
103'h387b4ee729604bea3000000000,
103'h0eecbd8056d10126f66000802b,
103'h2af4a2800e4c500e1e00000000,
103'h1a87b6ac1d390d8e7600000008,
103'h11007ede882db00e8469676802,
103'h30d992fb22b566baa200000000,
103'h2683a83eb4b5e5992a00000000,
103'h2b7a0d90648f78944c00000000,
103'h0ca980708a1320d3005dd079c5,
103'h3606a35f348d2e636400000000,
103'h05192d088236aed3ee00000001,
103'h04e19c4af93d52332400000000,
103'h2a398421bd567f3ba600000000,
103'h18a48ccb82381b869e00000000,
103'h3c9cc3d8ad719fa85d00000000,
103'h22cba9b9c5162c73de00000000,
103'h0337e1ce02b2f04c8a7e1ce020,
103'h1efa991de47e9a064e00000000,
103'h3cf56bf466b67bd45000000000,
103'h0661de7344b114f23600000001,
103'h14e47d6600a680e69c00000000,
103'h261a0ca547085f59e200000000,
103'h1cce35eadcecdcbfe200000000,
103'h3938db04c306e9652a00000000,
103'h1b549510ded51f5006f549510d,
103'h3e16d003970dfa54c800000000,
103'h28e16a5033628f65a600000000,
103'h2e98e15cb0795f693c00000000,
103'h375741ce585ac9b96e00000000,
103'h1ceac19006f3ab161e00000000,
103'h188c3ba67c4aece47600000000,
103'h089045229835ae747c52f5ab72,
103'h260dae07f0c1ea1af800000000,
103'h1ee5e0a6b8522f3d9000000000,
103'h1ab1be5ba15fdd45822c6f96e8,
103'h14c888f4fe45bdec3a00000000,
103'h24150202d8f77c47da00000000,
103'h2623652bacc0053cd800000000,
103'h2283f79212d5073fb200000000,
103'h3c44673df8f86c6b5f00000000,
103'h164a94d61a7c63fd7000000000,
103'h09483eb618c0cb3b6ac47ac6b9,
103'h2705edd2ee0b60118400000000,
103'h1898a42f76539ec79c00000000,
103'h0223c6f75c598c9a8a3c6f75c0,
103'h062b4dbcb4f230ca0000000001,
103'h24f39fbd7715f7c15e00000000,
103'h2ec751cfbe41457e1200000000,
103'h30eea2a9a334e53b8a00000000,
103'h0e6f801e10fc370b4836000500,
103'h20e28e5c80ead9b4ea00000000,
103'h2a6b945c4e5a59d2fa00000000,
103'h3335dfda313ce82f7d00000000,
103'h1c3510939aa87c8bca00000000,
103'h193078584ede5c65fa00000000,
103'h1416b9d1eb136cf99600000000,
103'h1e57551e8343e551e400000000,
103'h1ad4d89a965a9f23ce00d4d89a,
103'h30fad8a276b1f4425200000000,
103'h14ff35105086ccdce800000000,
103'h2316fe77c081a57f5e00000000,
103'h3572ad311480da8fae00000000,
103'h1e28fb0e3697d9076e00000000,
103'h3c913d2dac0a86388200000000,
103'h2c804c2a0b338146ba00000000,
103'h1af100a5c6c4be746600000f10,
103'h1ee28fb133450a9e7000000000,
103'h196bf7c40e360b443600000000,
103'h3effe60f6d189af56a00000000,
103'h2ec755a1848492b97800000000,
103'h255383a8028478c8e400000000,
103'h0f24bc4cf14bce6a6880462430,
103'h062c0036149f52126a00000001,
103'h2b4bdf14a4c40e5f5a00000000,
103'h12f050acaaf00e956e00000000,
103'h3d193b0d963bedaa1200000000,
103'h168df3d8e92c3e56be00000000,
103'h06a1feb6a74579645400000001,
103'h187a17f3bcd36d3d3c00000000,
103'h16423fc642756bf3e200000000,
103'h2b465542dcef83e7a000000000,
103'h2876a9163231c3ade200000000,
103'h0aec764dde7818f0be00000000,
103'h2b35b0c2c6eec206f200000000,
103'h0ef4572b90db3854d068080048,
103'h0ca2817bfd10e91796d974bfff,
103'h3e826f7a4a0540432700000000,
103'h0eda766956a7c1bf2241201481,
103'h25213f5f562a31396c00000000,
103'h0c4340aa2504a7a2c4a3f3d572,
103'h2f762b0c8b25e7021a00000000,
103'h1cae55b2166927ac3e00000000,
103'h208e4216c4df52b8c800000000,
103'h3a985fb4e08da86adf00000000,
103'h38a724f5c11bea81a400000000,
103'h02dbd138bab44a3684b7a27174,
103'h2179a527f55b6f2c4600000000,
103'h04f6cbcff63740650000000000,
103'h0a019ae2d6b0e58cf400000000,
103'h112854775ca7b15cea40518d39,
103'h1103584266a94c3fc22d060152,
103'h0739cb39b6d1a0b71e00000000,
103'h30a77e9606d4f8f98400000000,
103'h32c6177f4d0ec4333b00000000,
103'h108c61c57eb642c940eb0f7e1f,
103'h14fbf84b717c5a488e00000000,
103'h0f3d2f888308bc0e0c84160400,
103'h10535fbf1604b4597c2755b2cd,
103'h1f785428e641e3e1fe00000000,
103'h2b538b5bf69543a11600000000,
103'h26ab1cd7950d97c9fc00000000,
103'h270b6a613f612325f200000000,
103'h3c706c44650c3ffd8700000000,
103'h381752098b17aa5ec400000000,
103'h2a537b6fc68816a32800000000,
103'h309d3c9ffe9f68acb400000000,
103'h344820f628f2e41c7a00000000,
103'h1cff4549d89020bc7a00000000,
103'h10ce13fc4cd841b2a2fae924d5,
103'h0d24f951ead786fc7cfbfffeff,
103'h061b47543aa59af8c800000001,
103'h2804797306ca944ab200000000,
103'h247dcc4e4ce5db9eee00000000,
103'h2ecf60dc36ea5511f400000000,
103'h20f87c669b6821604200000000,
103'h0ec732e9c937823c7803811424,
103'h05607db7aa2ffea31200000001,
103'h06dfa42478f7318cdc00000001,
103'h3e491fa33d57af448600000000,
103'h101abc8242375368fef1b48ca2,
103'h2c23db9dc080730c3c00000000,
103'h335cf95c529b2f8e7f00000000,
103'h328d48a7bebf0b2c4100000000,
103'h2f154737b31c04889200000000,
103'h2cd49930a4a94d305000000000,
103'h2d145e35d2be94680200000000,
103'h3eef52c97e932d98a700000000,
103'h108952896ca78bce78f0e35d7a,
103'h123f56d1ea96de97f800000000,
103'h3a9ea84abb2031216500000000,
103'h32bc8e2b8e5f87f34f00000000,
103'h2b6da1a508fe303e0a00000000,
103'h0ec640ecfababe69984100344c,
103'h1eb5becce728600ea000000000,
103'h28c56dce34eea0fb9a00000000,
103'h0034a4c2d2a45fc8806c8245a9,
103'h20a20bf57b69cd96b600000000,
103'h3aca3191ba9e72598900000000,
103'h3c1ab73c9b407e4f0500000000,
103'h3359dde3160aafe0bf00000000,
103'h3b3d64521325671d5b00000000,
103'h3e8ab857c57f45007000000000,
103'h3e767eb6febca9528200000000,
103'h18a2c3653f4761aa4600000000,
103'h08d9b7f43cbde06144322bcabc,
103'h0b3613a09460a3c6824d84e825,
103'h1111b44d5c3a5bbabe6bac494f,
103'h14a9fe4ca6706f5b5200000000,
103'h1889a9f6368223a8ae00000000,
103'h162736010a2c21f55400000000,
103'h2a2565d262b5cbeb8a00000000,
103'h195df15e7add01ec9600000000,
103'h2f06ec45e40267bef800000000,
103'h38320ad5fc60591d7300000000,
103'h0e894b5b6a6745635600a0a1a1,
103'h089657cc64995039540783fa98,
103'h3a806629f2229b94bf00000000,
103'h126cdc467ab8f3612200000000,
103'h26b9ab807739598b1600000000,
103'h256dc01dc8a635d19000000000,
103'h08bb24f46e5fe152067262d334,
103'h1e2b255fd2cda16fce00000000,
103'h2e54192c5a88c6643c00000000,
103'h36b66683f8b3ebc41000000000,
103'h04bee9ad280804f06a00000000,
103'h03274e285ebe6b746450bc0000,
103'h125d5413637d55218c00000000,
103'h3c1c2062a4a4a349eb00000000,
103'h208ed875f601f75d4c00000000,
103'h2d099579b51e17bff200000000,
103'h1642bdf1d4acf035e800000000,
103'h24f93b8b82b685af9c00000000,
103'h16545c6f18f943a17200000000,
103'h3eb174affcf27f2cf400000000,
103'h1c2ca4b0d246db9c0c00000000,
103'h0f54c4e792f8504c0a28202201,
103'h03336acdee24f4fcdc59bdc000,
103'h0f0b5455bc79b9e46e04882216,
103'h18d5bd0a7ead24b25c00000000,
103'h36e7015b4cb879081800000000,
103'h24f095f8268e36129600000000,
103'h031f1f91dd75376de423b80000,
103'h1ac763100165cd660a031d8c40,
103'h321ccb408284ecf7e700000000,
103'h172aac791e4c5007e600000000,
103'h20c6c3c451691b486a00000000,
103'h06d8127d6693c7c18800000000,
103'h2d4f2e9c875a8b85d800000000,
103'h174b37b38d329e033e00000000,
103'h1e9390d27881cc9fc400000000,
103'h37450539d0cd04535000000000,
103'h348a4162ae609525c800000000,
103'h392a091166a59a5f9900000000,
103'h08fc6ec35b2fdbc248e9da8089,
103'h1350a1151559e4d3ae00000000,
103'h2a71d7ba1c5653970800000000,
103'h32f3a384eea6f4ac1d00000000,
103'h211b09af5b18cc663a00000000,
103'h2a724b9c0c0c6feb2800000000,
103'h0723725c6e27799a8200000000,
103'h012aecb3d899c53690e258f534,
103'h2ad95bb75ebd3792fe00000000,
103'h2ca0972120e82446d600000000,
103'h3d7442760ac17ffe3400000000,
103'h3a6f67657662171f5500000000,
103'h1104518b74d659955e16fbfb0b,
103'h065673446f45c0fad600000001,
103'h1a90b944414a12864a0242e511,
103'h3a8c7f4246a085cab800000000,
103'h10ea5c5fa0313f0ef85c8ea854,
103'h1a1e93125abdbe513e00000000,
103'h12988abfeaa81ab0e000000000,
103'h0c5c94f3c4c6adc33a6f5ef9ff,
103'h0ac124f2595f38832600000c12,
103'h2b56f3ffe4bbcd76ea00000000,
103'h26aa815eae7cf2694200000000,
103'h0ca6296e5ad3e669267bf7b7bf,
103'h37687f41417e67c7d600000000,
103'h3a8a0d974d2491363100000000,
103'h20676964428d10777000000000,
103'h36c1b79a7d171e0ebc00000000,
103'h26efec39de7e8772fe00000000,
103'h169c88a115403f0d7c00000000,
103'h136db63e7d302b475a00000000,
103'h12cbf45352ccb3e86e00000000,
103'h0f415076e63a6a26ea00201371,
103'h2935340d79065e7a3e00000000,
103'h176956b18747aef12400000000,
103'h02cda49cef7ce2fe9c939dc000,
103'h00fea670c4e639b022f2701073,
103'h246a126b86b3de4d1000000000,
103'h00dbdce086b284bdd4c730cf2d,
103'h22955646ab1c97295c00000000,
103'h32cbb2ab6af87409e300000000,
103'h06e848c04c8dca508e00000000,
103'h22b8bd223e597cfbf800000000,
103'h073bb6420741c5bc4600000001,
103'h14db468b28fa82de8400000000,
103'h0c734ade2e3639208a3bbdff57,
103'h12991981c3117fabb400000000,
103'h191865215084ca89e200000000,
103'h22d9767d231de40ba600000000,
103'h16950ab77b36492cf600000000,
103'h3a86d8125e0fbfaa1900000000,
103'h208a2518f4a4ca619400000000,
103'h16123ca96f2ba273f200000000,
103'h2eb838458eb5c78ce600000000,
103'h02947d0ea4c8043656f43a9000,
103'h34808181d4803c7be400000000,
103'h1c1150569714b98a8a00000000,
103'h32cdc19f4c953b0c5f00000000,
103'h173ffa74e8a68b62f400000000,
103'h217a3780da744d024000000000,
103'h3e34b108b0b447772800000000,
103'h3503e41b122e7ef80200000000,
103'h34685239d1633000b400000000,
103'h1e734bbb8567141bc600000000,
103'h20f2923f7acf66559600000000,
103'h1526203a9942b2111c00000000,
103'h1a882d2db935445096000882d2,
103'h334d6a218f5b648b2f00000000,
103'h0e79bb3128e391b8e630c89810,
103'h247572965a30fbda7400000000,
103'h12b3dc0ca8aab70b9e00000000,
103'h382789d38c2029a1f800000000,
103'h2ef69c259ed405aea200000000,
103'h0ca9403098fb8f822e7de7d95f,
103'h048ce01606f22ba7ce00000001,
103'h271b3707129b6bd86600000000,
103'h16c9b79a17284bee6c00000000,
103'h254c3ddbbf4382f57e00000000,
103'h0aca539f940d3a8f9400194a73,
103'h373a950b3859786b5200000000,
103'h3546424f4223cc0ae600000000,
103'h097a3b81b85e61161e922d4bd3,
103'h1cf1b7a9aca4a3656000000000,
103'h02766e61341edee7187309a000,
103'h22549d8410109690c400000000,
103'h035698b1d48704f1fa40000000,
103'h1cb6f4f5b6dba2760a00000000,
103'h20bbf49ef8323b27de00000000,
103'h1adfd32f54e9301d94001bfa65,
103'h2714485076a524bc8e00000000,
103'h04cfc2639084f7ebe200000000,
103'h1a66deecb699403c58000336f7,
103'h2930369dbd69029fea00000000,
103'h0ae2be6c56cfe18ca00000715f,
103'h253a6af77e00182a5c00000000,
103'h0e170f6e88e2d696b201030340,
103'h2e8cf421ec1d418e3000000000,
103'h0c6bdb753b3450fcbabfedfedd,
103'h3f1aa4552ac1451ea700000000,
103'h30c9855f772d2093e200000000,
103'h2a5b3d007547c4e90c00000000,
103'h100a362fa5114a48827c75f391,
103'h32ed805b8e6c8748f700000000,
103'h3e920fa62176bd789c00000000,
103'h0063bf8492643dd42a63feac5e,
103'h397d344c12f64d7a4b00000000,
103'h14a7f35c135a0cfede00000000,
103'h3e3f39b50ad7414af000000000,
103'h0a4d3d869e7f34a702134f61a7,
103'h28bf7f2c5ebe6e5c0e00000000,
103'h19280e4c680babe2ac00000000,
103'h1aeaaa6b50cb2b0f0a03aaa9ad,
103'h288487d528f3395b7200000000,
103'h169d99e602dde3c6c200000000,
103'h21751a52ec626b9bea00000000,
103'h155846a283000581ee00000000,
103'h16069e0123751fd4da00000000,
103'h02a82ebb36cd66775cd766c000,
103'h3127a33c0ed404787e00000000,
103'h0b098358d17c3333b600000010,
103'h26eb68f780a3d66fc400000000,
103'h25426e6b0aad59c89400000000,
103'h1b66da55f098c2c014ffecdb4a,
103'h1e5f4ab954db312b1e00000000,
103'h32d3ee5071420b810f00000000,
103'h06ec68574ea1563a6200000000,
103'h24b23c26c275448ad200000000,
103'h3210d2b64961ace22300000000,
103'h174a9a70ef13e908e400000000,
103'h28c66daca024bbbf2c00000000,
103'h0ae39722b66f56301a00038e5c,
103'h2f760523a135c3dcbc00000000,
103'h1c6a2006aa195aff7200000000,
103'h377223f29a8f60231200000000,
103'h329ee39db6f98029bf00000000,
103'h263af978ed6ba41c5800000000,
103'h390cd330e10a87ba0e00000000,
103'h36f807e846458132fa00000000,
103'h0e729cc2be525463da290a214d,
103'h1ce6b1c6f64a5c4c2000000000,
103'h18c66ae784bcf90ee000000000,
103'h32b0abc222a3aad5d700000000,
103'h14e06dcfba6a15bd5a00000000,
103'h346284412c1ac17f7c00000000,
103'h0a2ef6fec0fb2f4f3600000002,
103'h24b862cb355db3906400000000,
103'h22e5796d7e8caa8f2400000000,
103'h197ca5cd25450d5a5a00000000,
103'h3d2e93ac462a86c7d800000000,
103'h22dbb0da9ea72c94fc00000000,
103'h3ce681995cd5c0414200000000,
103'h157dfce73eb1711be200000000,
103'h135a858f7a97f2b53e00000000,
103'h146194ff8f15ef9c7c00000000,
103'h360fd104a170752bf600000000,
103'h3493cd4af6d20a2b8400000000,
103'h30c93aad2ce1db302600000000,
103'h26969ac4a375a87b1c00000000,
103'h2c79ea78923ee3284800000000,
103'h12cdaf587ad57decea00000000,
103'h2ef37e63e74f68657e00000000,
103'h36fb289f791d17bdf800000000,
103'h23787b5627109621de00000000,
103'h2034b1351d0bbec15600000000,
103'h18c66500fe843a177c00000000,
103'h36a781325eb8eb4c9800000000,
103'h0ca5b521b77f504d98fffab6df,
103'h08b47f32ec26d17ff64957268d,
103'h20cf080578cc86a1ae00000000,
103'h386dcaef808105d49b00000000,
103'h30c5792623500dda1400000000,
103'h1e9c77aa5abdd8c99400000000,
103'h389a47ae8a8351efb600000000,
103'h0c649e54691fc99a12bfefef3d,
103'h22affacee2ba11489c00000000,
103'h184b65236f1eaf9d0600000000,
103'h2aa4a84190ceaa6be800000000,
103'h08813d4f6a1a0f8f564d99601e,
103'h0e7d9bf754beb7d0e81e49e820,
103'h36340be7dd3ff5205200000000,
103'h0c092b756abd9117a65eddbbf7,
103'h34acf56ee0f19cff8400000000,
103'h076acef7aefac874ee00000000,
103'h2ee7605162a7bde3d000000000,
103'h32a3e6cb6b128cdb7f00000000,
103'h211dfe5d18f9ed2ce000000000,
103'h3089b2ee4a9dd3f84a00000000,
103'h2ef02ff46abbd2556200000000,
103'h10fe6ade5c458543ac5c72cd58,
103'h1a1f32a3cb35b538180000f995,
103'h3e39e7961b3420167400000000,
103'h2af27080b65352ba3e00000000,
103'h0366cbc0b48d3a505abc0b4000,
103'h3620ac445f7faad11000000000,
103'h3710420022e67691c400000000,
103'h1033f7d2580722d622166a7e1b,
103'h20ab005ece1764d64400000000,
103'h24af433b9f4b5ca89e00000000,
103'h063330e97ef65d076c00000001,
103'h0c9d952922a5a0430c5edab597,
103'h2b0f1c3eead8d12c8a00000000,
103'h1698082af7766655ae00000000,
103'h236c50bfa08582949800000000,
103'h2e36f65bb71d8abf8e00000000,
103'h1ca73c3ada89db7f2e00000000,
103'h34f0534688c0d1dae400000000,
103'h02afd0a7e4680e15be00000000,
103'h30f4d09dd858615c4600000000,
103'h15575b535a0832042a00000000,
103'h1543c1880afd02a20200000000,
103'h1af0f9979e545df55c0001e1f3,
103'h06063fbcf2981f7d6600000001,
103'h0973e73e8e89191506fd7f15c4,
103'h26e9c0c4548f58d1f800000000,
103'h0c5c9cec1c034010862fee7e4f,
103'h1223d70942ed00d4da00000000,
103'h0c8330a3d1499dc0f8e5def1fc,
103'h126ba353626d74ca3a00000000,
103'h2ee36ed4eef0a56e0a00000000,
103'h275e7a67035c48c16e00000000,
103'h20c686cdf03fb7965c00000000,
103'h2d7830f5d69e31fd5e00000000,
103'h1a974fe7f664b8cb4e00974fe7,
103'h36a7144822dce9c12400000000,
103'h16132169bd7439a91c00000000,
103'h24bee621b41b4df13e00000000,
103'h0b08dcd70b2e6f5afc00000002,
103'h26b78c57aeed557cb000000000,
103'h2443259978f63253ba00000000,
103'h2042f8845eadbeab6800000000,
103'h115e196084f0e444e2369a8dd1,
103'h0aa7a997a433dcc94053d4cbd2,
103'h34de8f4b7691f629c400000000,
103'h160ba75301399fc16a00000000,
103'h16e67e05f5182f0ce000000000,
103'h1cb238fdca23d65fe000000000,
103'h06b1d0bee30a5465d600000001,
103'h27435ea9bebc8d63a000000000,
103'h070e8c56046e5e228200000000,
103'h1cf1e90f2ab1bccc4000000000,
103'h3ef91c2830c049224500000000,
103'h010aa3a70eb232316ede6aec3e,
103'h02d8b8898cab4e59a044c60000,
103'h06152b8e8cb5f200ae00000001,
103'h36035b5fce8eaa8a3a00000000,
103'h16b1d45356a3d618c600000000,
103'h05127f784ca731789600000001,
103'h3f1e78f6e35905cbec00000000,
103'h04e06476276b85443800000000,
103'h1b30fa7fa489fe3b1afffcc3e9,
103'h062566a1e96a62b14000000001,
103'h3ec1043cc49b5d30e500000000,
103'h18b5a7a38ac0c3d2cc00000000,
103'h1915d04e8a81c80f9000000000,
103'h3cfff734a3376fb31d00000000,
103'h0b5480cbfd4d4001a600001548,
103'h1a446794384d37364802233ca1,
103'h36f5122f42a1b8024400000000,
103'h1d2784d9dee61f967e00000000,
103'h2691673794db31c5c000000000,
103'h2b488996f202b69f9e00000000,
103'h294ce32c98941dd73400000000,
103'h2af2f4c482dca76e2600000000,
103'h097f25f2ed298a9abe2b57b429,
103'h3ce688e7161c7f5f4000000000,
103'h2250a27ade9ba5522c00000000,
103'h214ed9e5dc822e394200000000,
103'h2229b8befed2d0b42200000000,
103'h0f2e2232e121aa99fe90110870,
103'h134f0b06024b6358fc00000000,
103'h340b992b5079858bdc00000000,
103'h324a5589e2c89091df00000000,
103'h2e5be29c96d429bd3000000000,
103'h0c8f1a49481e7f47124fbfa7ad,
103'h2b0db54ef97a61e3aa00000000,
103'h1b05d5e084097c2cf2ffffffc1,
103'h2ec68703ee17317bea00000000,
103'h195b61e48a1d075c6e00000000,
103'h0b0ebc0c38e38e605e00010ebc,
103'h373c7817913ef044e800000000,
103'h2473b04fdb4dac512000000000,
103'h02c21a04108a2468b008000000,
103'h2b2d8b14b6fdd4b88a00000000,
103'h0a7c8a85b8bfeebc9c0000f915,
103'h3b0a7a3ba4ed79d15200000000,
103'h06e61642ae6a04570a00000000,
103'h234bd6b26a747e92ae00000000,
103'h34af6bdab15a94d55e00000000,
103'h3ed2efbf92a66b87c900000000,
103'h2ee3ed75c755d7627800000000,
103'h0c5eef830528c7220abf77d187,
103'h144e7022f30cb497d000000000,
103'h0c9885983e6ba41ad47dd2cd7f,
103'h1689069552ba143dc800000000,
103'h26cf5ef4de5299d60600000000,
103'h3a3e7e7674dba06b5a00000000,
103'h02ba528fdaaaff6038d0000000,
103'h0aa1cac416e97dd6ae000000a1,
103'h2443573618a3d0668800000000,
103'h1c377d7e22459b2a9e00000000,
103'h0a0744318688f260b800000000,
103'h14820a4524c06fdeda00000000,
103'h32e64e2f6ec7b4106300000000,
103'h2aee62804349be558600000000,
103'h073c11fbb6300c84f400000000,
103'h2812b3d7e11e6f053800000000,
103'h2ea9c592e75a8100ee00000000,
103'h22088b5e4e6d34d8ce00000000,
103'h1ab10f7f3d16fa6bb60000000b,
103'h0889a025201f85ca044b12f792,
103'h18809fd03ad095494200000000,
103'h0ed2207c455a356e6229103620,
103'h1290d6011cdad53e9c00000000,
103'h156685f1aaacf5bae000000000,
103'h365bbbac3c3dcbbbfc00000000,
103'h152186b012a451ada600000000,
103'h3441872249000d59e400000000,
103'h323c5cd31d219409f700000000,
103'h18e4283ed2631b2c3e00000000,
103'h3cc9bf66849f77ff5c00000000,
103'h3253a83bdc83a03e2f00000000,
103'h32dd9e6b1b4d5fa4b300000000,
103'h0e8928a44ca107e08e40805006,
103'h3c97ce09be7ea64ba800000000,
103'h2e45eb6e8d07ceeff600000000,
103'h3c77a911889f9cf9b500000000,
103'h26f6c65936e588684200000000,
103'h1d16eb81745d3179ca00000000,
103'h10b5b6f55b53f7d302b0df912c,
103'h135c5159376ae3547600000000,
103'h1ea288b6c7209a49d000000000,
103'h20ce487c9b7ceba30600000000,
103'h175739bc381f7459cc00000000,
103'h273422ced8edbcd66600000000,
103'h2d7bef35ee44f6929e00000000,
103'h38e455e6d47919617600000000,
103'h20c9a83ac0f508976400000000,
103'h3ece6ee878d95e7e3800000000,
103'h36c0f26c98a306b8f800000000,
103'h1af86c83597175a1720000003e,
103'h14a8fffb8e32680e0a00000000,
103'h0c4e9c0b282ad49162376e4db5,
103'h3ecd9698fcd3d48cf000000000,
103'h0aef97dfcb2270981a0003be5f,
103'h2c830ec808f007311600000000,
103'h1e48edbe52df9f10e000000000,
103'h3939a1460162add8eb00000000,
103'h0efe295a9eab9b973c5504890e,
103'h30e5220756e53cdd3c00000000,
103'h1abc21e524e36637da0002f087,
103'h1672c0d3d4c8883f3000000000,
103'h148c0d9b6e84aa245600000000,
103'h2f50f5fa46f76af82a00000000,
103'h20fb1b365a8378939a00000000,
103'h3688a6aa48d46e8de000000000,
103'h20deba5d68cf89c43a00000000,
103'h3ab97834de58306e8300000000,
103'h1a8ba1048136eacbec00000117,
103'h14e14267baf06300ca00000000,
103'h190b5258d67c04054a00000000,
103'h0404ec0e2b5d466d0600000000,
103'h0e56b632036898c5dc20480000,
103'h1adf6b21c66d84d4060df6b21c,
103'h2158831256c43b060a00000000,
103'h3d4d9f0830a3a627d000000000,
103'h02a0016b10fc293a26ac400000,
103'h0d5afc93cc49c84256adfe69ef,
103'h1e837c908ee9c9ad6600000000,
103'h057037935c44c6413200000001,
103'h1d0098bdfac842d1c200000000,
103'h028d2322bf387a651ec8af8000,
103'h366375c9db3913231800000000,
103'h3923921e5ec63645d700000000,
103'h172874b41529ac0fb200000000,
103'h2ef59a1b8d4d3e2e1000000000,
103'h04fb39e82375b2e22400000000,
103'h3739ecd7d16b4cfdb000000000,
103'h063ed60d556686e5d200000001,
103'h2b6d6b528ca073bda200000000,
103'h1ae93ec5d2df49caf60000000e,
103'h2cdac51b3e4cb51d8200000000,
103'h0e37986e5935f3e3561ac83128,
103'h06faf2a74710b8fe9400000001,
103'h085ec09dd448516cec0b48f89c,
103'h1ea1d85f5a4344143200000000,
103'h3331a53e64a204b20900000000,
103'h20f76600c243dd116200000000,
103'h12cddfc1b675824fc600000000,
103'h1aecaaef976ce8508a03b2abbe,
103'h3e4eba31a93ac8124000000000,
103'h0552ce25c5277301d600000000,
103'h0e9abf2b42762d337e091691a1,
103'h0e58328086c8fb594224190001,
103'h24828e265663ba848400000000,
103'h24e7b1de64bbed050c00000000,
103'h277448984b3e7b2b6200000000,
103'h2d770c85ae262d09c600000000,
103'h3842cbcc549a75a21100000000,
103'h1a72459780118227be00000000,
103'h205dac67b9544df41400000000,
103'h32878e6352c6938b9500000000,
103'h30d79d68b5243ff34e00000000,
103'h04c2221026abce56a000000000,
103'h1abe28df56836bbf540017c51b,
103'h290e7da29c458dcf7a00000000,
103'h092565f17703b6aed21369afd2,
103'h1f608e339f1234516e00000000,
103'h184784cc67379a42e400000000,
103'h2ab1e724849828768200000000,
103'h1961d74c1edfad42e800000000,
103'h3c157e22889194676f00000000,
103'h3edb594a62f36bb38c00000000,
103'h28d8ceb51e08e9d61400000000,
103'h176e6c965ee443207600000000,
103'h22e3b7ba86bd11d59600000000,
103'h36ea97461d2b7e6bf400000000,
103'h2ee4e2853f0f36267a00000000,
103'h04e8179a74f9cd6c9600000001,
103'h38cf8fd022deaff1d500000000,
103'h327419db66c6c78c4900000000,
103'h084422529e96575c6c693a8779,
103'h1c2360f0500a7137d200000000,
103'h24fc6cfa994e938a7200000000,
103'h10b428f6b471f47ac2211a3df9,
103'h2532ac7f1b6e61755c00000000,
103'h16478763ea228a6c1000000000,
103'h1866d3808e5536eb2a00000000,
103'h34d4b327a49cbe4f1600000000,
103'h06b487497e0391cfa400000000,
103'h3002bce0b2d844f74a00000000,
103'h06737ce3f88ccc40c800000001,
103'h2d3973d26a8f89217a00000000,
103'h369c290ff10306057400000000,
103'h3e02701d1d3c79d7de00000000,
103'h3840fc2192d8a2e7cf00000000,
103'h2c0c5466d0db1304ec00000000,
103'h0b6735cd8a1c0f267e00000001,
103'h1ac51d39b728638d5000628e9c,
103'h075f7e7dc28f995ada00000000,
103'h04d282a99c54b6949000000000,
103'h152099da62b435125200000000,
103'h2e8ac031a686b7bbee00000000,
103'h011d4a163ca7519650e24dd646,
103'h123f6d55ab3211c7f800000000,
103'h02b64729ab4f5bde3454000000,
103'h12e1560ffe8ec933de00000000,
103'h0a931cb24145105d8a024c72c9,
103'h3eec34ead326666d8800000000,
103'h1f775eeb5eb9831fc800000000,
103'h2851e4ca1ca5b80a9a00000000,
103'h30bb33dcba1d16f5f800000000,
103'h3869934ce36efbc01600000000,
103'h123e592a922a2f9cd000000000,
103'h0ccca2280a93c2e9b46ff174df,
103'h2300a3301ed21c144600000000,
103'h3351bb2e2a9ebe3c5300000000,
103'h2711ceec4c9f616c7000000000,
103'h2efc12473ef11c9a9a00000000,
103'h017a188be702eb86e63e820966,
103'h30ca3ae4d4fefdce2400000000,
103'h0ab91b7a1479165a0a02e46de8,
103'h31475d7bc443513ede00000000,
103'h14c6bc180efc6cb8f200000000,
103'h2149063b3e43ca34b600000000,
103'h3eca4e2c920a864cc500000000,
103'h32c4ac77f2538c880300000000,
103'h29025c02331ddab49600000000,
103'h2f3c784564e2872c8800000000,
103'h30ba5ebd4ce4e32eba00000000,
103'h0642cb81fa215b741e00000000,
103'h111ec4ceacdbba316c21854ea0,
103'h0a1898cff21e85b36600000189,
103'h2af4f3fdc23d4a821200000000,
103'h16b6325a4f55e3520600000000,
103'h3c98cc2af84ad74fc800000000,
103'h1157202d0e0109aa16ab0b417c,
103'h1633f9e28a99d5d50e00000000,
103'h1e4e1e1a1af0f6021c00000000,
103'h36be25a3b124efe4a800000000,
103'h0579047d10730dfec200000001,
103'h2334ed00873133a27400000000,
103'h0a8aab590aaa381f8411556b21,
103'h0cd15fb3acdf25200a6fbfd9d7,
103'h003d03f2f669d07914536a3605,
103'h051bb631053b302cc200000001,
103'h0e2b9c118478341fb8140a08c0,
103'h24e5ba118a93ea50bc00000000,
103'h267efd3198bf86624200000000,
103'h1e8210cabca54073cc00000000,
103'h1cc05490a2243da56400000000,
103'h1f76cc7642a64e702200000000,
103'h2ac12eac9e66a300c400000000,
103'h0ecb17453cdd6f77066483a282,
103'h317a4051a69e9e23a400000000,
103'h364da7037469b568e000000000,
103'h3cc75c2566e3f5ba8700000000,
103'h22a7b4481d319cbdfc00000000,
103'h02657be1d8f8f8e362e1d80000,
103'h0ac1e19f3aa0ad2b7e00000000,
103'h0687fcc57e06290d5600000000,
103'h29320da648c80aac9200000000,
103'h270dbb450f5007721000000000,
103'h3ce261c7368215185800000000,
103'h0f57b574dc8fd05d6603c82a22,
103'h1ed3322fd97232249c00000000,
103'h3716b99768c9e7997800000000,
103'h1caa4871069d19c95000000000,
103'h38bfec62feb3d360b800000000,
103'h306560b25b5e1bd1c000000000,
103'h037d0726551e0834be00000000,
103'h3a5e9533c48368e71800000000,
103'h3add3d0a8600700d6d00000000,
103'h390fb842035f05413300000000,
103'h12a04f4b3c3c424bb800000000,
103'h3f4eee89364bfa8dbb00000000,
103'h3080f6ae48ec49d8f800000000,
103'h2ab36ee0c73b38622e00000000,
103'h2544ec5478bc2f107600000000,
103'h1d12ac13e26f9df13c00000000,
103'h0a2c666106b48a45b400000005,
103'h01326a8724c7365996fcd0705d,
103'h3e73a70f6ef39cba9e00000000,
103'h337112a831260741c300000000,
103'h0ade1c322e99ae51300000006f,
103'h28ffb001e00ac0f96000000000,
103'h2ae87a2b2ae8dd2b8e00000000,
103'h1ac4e10f12e88d2d7000000062,
103'h3cc74f34bcd107589b00000000,
103'h0b636bab9895e867ae00000163,
103'h3b0a491bd45d379c6a00000000,
103'h169a03b79ec0a3480200000000,
103'h05124b80dacaec63d600000001,
103'h2f5b9aa2b164f01b7600000000,
103'h333ad22c35773b9c5100000000,
103'h0877415222d2d63f0052cbb691,
103'h3e7453c0150da86b3400000000,
103'h0f3c5291de84e9bd56022048ab,
103'h0e69417f1cf93d7d6c3480be86,
103'h030d6c08ad35900f4ad6c08ac0,
103'h1a846cd13a9ed18e6600000846,
103'h07091604feac3d971200000000,
103'h1112a8f61930aa684ef0ff46e5,
103'h371579649f39c06d4c00000000,
103'h0b4dd9e26f4c696364000029bb,
103'h18250beea561e2c80200000000,
103'h24a87b91eeafbcaa7000000000,
103'h085c959d86d4c89914442e8249,
103'h0a4a70166b7d442b04094e02cd,
103'h3a84b3f2b2d9d9c88a00000000,
103'h0e20da96fd2449def610244b7a,
103'h126cbde5b6a8fdd1a800000000,
103'h1e8d69cd86c9d868a600000000,
103'h142b59e05836964e5c00000000,
103'h3ca323bbb6c4001be300000000,
103'h223f37760aef59fc3c00000000,
103'h0084490208927db7f28b635cfd,
103'h229332f6aad1b52dfe00000000,
103'h1ed8b339ab55fe300600000000,
103'h12e233988ee93126b000000000,
103'h10db0df3acc1e4605c0c94c9a8,
103'h16666606bea417f8ea00000000,
103'h06c37347ce7f25ec9600000000,
103'h22767eb8e4e58bf35600000000,
103'h0d12bb50aca8ff3b24dd7fbdd6,
103'h2470dc48cf1f7df40a00000000,
103'h3b731539dd323944b700000000,
103'h1ef4741780a3158d8400000000,
103'h295b5ee87a162ac76000000000,
103'h1e6b48f4980a9edee000000000,
103'h249ab0f4c265fdc75a00000000,
103'h04fc5239a0d146bbf400000000,
103'h2601090c056bf7b0b600000000,
103'h011beaa5ca6849ea56c21a4810,
103'h35416b1e716952f65c00000000,
103'h2acce95e70853d9c2600000000,
103'h0329ae5a66c6a8ba96b9699800,
103'h1ef26b07109392190600000000,
103'h0423719e12bd40736c00000001,
103'h1abdcb2b70afab7a7e00000000,
103'h20dd6254f4d31d189000000000,
103'h0ec3a2390e90e8440240500001,
103'h0d3d7436306e4a98f6bfbf5f7b,
103'h1d7486a6bf31ecd20600000000,
103'h1f5b4491cb6f61083600000000,
103'h16151f9566e3e7aef400000000,
103'h1d5fe2dd073f2c40be00000000,
103'h1318f0bd9c544bd62400000000,
103'h0703eb7038b42eb32a00000000,
103'h055e472b0acd1f70c600000001,
103'h289c8a94d0d10ae0fe00000000,
103'h1519fa3f542f520c0800000000,
103'h1aebb5bffccbdca0d800075dad,
103'h1a719ff3d0e5d6e02c000000e3,
103'h22c4a9986cd18ca02a00000000,
103'h3ce8be1e06432c93fa00000000,
103'h283c24afa807d62c6600000000,
103'h125b67e224f0944a6c00000000,
103'h0f6081f4cf2cb8fa1690407803,
103'h343728a7a08820dc3a00000000,
103'h2250fbee6ee8a2d10800000000,
103'h3972a561a51fcb78aa00000000,
103'h3284e31f4670c7671900000000,
103'h3cc3d9d6fee36cc8bd00000000,
103'h268af16af0684fe80200000000,
103'h3e3aabcfec2c29bf0100000000,
103'h3c0a31ad92b71b29f300000000,
103'h3f4a7ef252f1c6f9df00000000,
103'h016e38ffcefbf8a7723518d3a0,
103'h32fa42f54d467799c500000000,
103'h10b276a9ccb4b09992fee3081d,
103'h0221c5883eaef38ede620f8000,
103'h0682db6091616a38ac00000001,
103'h18dfe9e052832fc0ea00000000,
103'h38836ff9da060b217a00000000,
103'h24dba6acf2e5f501ce00000000,
103'h0ee2d0eeeb6964fba830207554,
103'h0a4b65698e450ba89a00012d95,
103'h193729a51f27dc978600000000,
103'h0128f9022873420114ce1d819e,
103'h1b00bd6100aa6ba632ffffffc0,
103'h2141e6bb80d364a85a00000000,
103'h36c81bbe9ad422095a00000000,
103'h29762d593c1608c4da00000000,
103'h049780f4f2de24837600000001,
103'h1e634036db5451dcb200000000,
103'h3a0264211eebd2d1a400000000,
103'h3175aa14be4f13087e00000000,
103'h22fef8cd395177299e00000000,
103'h07666c0928c7213e5c00000000,
103'h05223121cac61a0b9400000001,
103'h22c9c90c112c8614bc00000000,
103'h3ec073fed54eb7368600000000,
103'h1308961b391880429600000000,
103'h0e17d975f6d8f4416a086820b1,
103'h14ed36dc4ae18a5ca200000000,
103'h2aef1a5758f963d29a00000000,
103'h173fb508eee69aaee400000000,
103'h38a8cffd18d5b5063d00000000,
103'h12eadf32ae156a0f2a00000000,
103'h370e78c4e8be3a0c4400000000,
103'h342b7629baa9193ef200000000,
103'h1f2f0e3d72b79203da00000000,
103'h23085b5766e3082d9600000000,
103'h16f712808512166b0800000000,
103'h30a403b5e91a71c26e00000000,
103'h06fa0e2a3e118442f200000000,
103'h0e07aaa26eb587f8da02c15025,
103'h3cf84f4836af96231800000000,
103'h30fb0a5904b740c58800000000,
103'h0b18372c42af900dbe00000001,
103'h2546e84272aa9a66c200000000,
103'h2c2b21517cc2d1930400000000,
103'h2abef083a009b9d57600000000,
103'h2c0a007b4d34db26f400000000,
103'h3204a080b6f3cbaa9500000000,
103'h28a9daece4fdcc25e200000000,
103'h1d11e6ec16026ca69800000000,
103'h3283acc0beac47937d00000000,
103'h152a4dbc5cbe2e7f9200000000,
103'h2cc4ba628f41db405200000000,
103'h2b5cf32ea36c28fcae00000000,
103'h3cf798a14f30e35f3d00000000,
103'h0e3e85a7788dd68dde064242ac,
103'h3d43a12d36856f2f2c00000000,
103'h388a97f344c3f4d6a700000000,
103'h173db7b603079603dc00000000,
103'h0421bad7fa922df72000000001,
103'h2a939487d2cfe5ad2200000000,
103'h068add66d6f1a0851e00000001,
103'h27461b1c8085350cf000000000,
103'h0b08eed607101273c6108eed60,
103'h285df086ad562d904600000000,
103'h1882d7e4775f1c664c00000000,
103'h1e995fc75ebd0cecf800000000,
103'h24351cb7373fe4d17000000000,
103'h30e0ec1ad4d94498ce00000000,
103'h28e2e90eb90e61500600000000,
103'h18440268e8ef4d6ada00000000,
103'h296228b012d236799400000000,
103'h2ec033c8aa1638e27c00000000,
103'h08f7837a127861928e47f1744e,
103'h1c3d347b8138955b3a00000000,
103'h1b7232e7ca3018d54cfee465cf,
103'h287967cda76d4d50ce00000000,
103'h2296d59600df80389800000000,
103'h312ca4f0ea58e8063e00000000,
103'h3efb09a70cefbd9c4100000000,
103'h16f987327d1c628d2a00000000,
103'h1465520eba176c343600000000,
103'h14b09d239110f366b400000000,
103'h3f54d03ea67645756f00000000,
103'h36e8c0f5fb26e2990000000000,
103'h2a99143a7b7bb2d7a600000000,
103'h1960d3b3306473cda000000000,
103'h193986929afd88081a00000000,
103'h3e887ee7725e5bbb4b00000000,
103'h20fe59d54c97e24de400000000,
103'h3aefe79acb2061355900000000,
103'h0645e92deb1ebb0aa400000001,
103'h2a9972c9260ea2a56e00000000,
103'h034b581fad548bd35a81fac000,
103'h26951fc416edfe9c8000000000,
103'h16ff489ddb3956bc2c00000000,
103'h30882c8240ce76804200000000,
103'h301fb30c16cdbf1e1c00000000,
103'h1c0bc5694755eba05e00000000,
103'h1ee5d662f6759eac7400000000,
103'h3cf93e18d2816415bc00000000,
103'h1adb1c4ef2673a78b200000036,
103'h0e8ab9a32f60789186001c4083,
103'h0a904297c93b94e07800000004,
103'h3e0b6a38d6c64e83a600000000,
103'h0507f5efa356911b6e00000001,
103'h3d6bbc1f2061fb544400000000,
103'h232ffae02469f143e600000000,
103'h112fce81a0d5ad63062d108f4d,
103'h14f5f0a6c205a8432a00000000,
103'h3d12a3e7523576c4ca00000000,
103'h0291527c262b676b8c2a4f84c0,
103'h2e79f254e23e0b52de00000000,
103'h39383f90a6cf5dcf0700000000,
103'h06fc350f94495023e800000000,
103'h24f5a1534c818fb48e00000000,
103'h2a1a7502927dc4c42200000000,
103'h157d5404b97366177000000000,
103'h22af90d5e28ddb1a0200000000,
103'h062b1dcaf60b2f1eba00000000,
103'h37283a749ababff49e00000000,
103'h38a31be260e5ddbf9500000000,
103'h34916367960e18342e00000000,
103'h120d8606ceb134168e00000000,
103'h2694d7c4c242977e2400000000,
103'h16d6e97755501d84f400000000,
103'h24fed8e97ce4f549b600000000,
103'h0b34e08fd2bbdec10c0269c11f,
103'h3e1c1c4cb6bab7aa8800000000,
103'h3445ef87c0ef983a5a00000000,
103'h00bfe047be0bb4871065ca6767,
103'h091ec6517551a40ed227b12fd3,
103'h22398b1c341184569000000000,
103'h350f07917e304aa80400000000,
103'h06d41c412169d5c43a00000001,
103'h16a4e577d578dd55b800000000,
103'h1cc752bd5a4cf996d800000000,
103'h16fb445972f1df0eae00000000,
103'h0f5f809d8eb931cc080c804604,
103'h272d92a5e4b476257a00000000,
103'h15748203f213f6c30800000000,
103'h1e086af8d8418968ec00000000,
103'h188e32fc6eb60b6cde00000000,
103'h22cd2ccc0cbe7665b800000000,
103'h0ec09cc1254ca9622620442012,
103'h2ec803794719d62e3200000000,
103'h2710f39a56da72ef5600000000,
103'h0d0fef2844a276689ed7ffb46f,
103'h3ecd611beab36a02f500000000,
103'h14d77c71b6c3592b3800000000,
103'h32fb6df5b490ba472300000000,
103'h26f9d269096836b8d800000000,
103'h1e9aad44fd63a4ae8c00000000,
103'h00eef223e25d771794a6349dbb,
103'h1906902e02f8245c9000000000,
103'h24aee87f42e716807400000000,
103'h3abf77895ceda6ae7600000000,
103'h0a33ab42009c8f2db800000001,
103'h3e0556123a5c06b71400000000,
103'h34cf253f068fb1f91600000000,
103'h2e800aec4495080b5000000000,
103'h031e9747fa642d4a565d1fe800,
103'h1959b2d168e438369c00000000,
103'h2af0d511eb02cf7e9600000000,
103'h0117a94b855c824ffe3a15cdc1,
103'h1cd385906e4d5761e800000000,
103'h32f38f1fae6500ad6d00000000,
103'h30f7d0e58c38863dda00000000,
103'h1afee229ff2c155d8a03fb88a7,
103'h076275be7123e6431600000000,
103'h231360b4ca22c86d1400000000,
103'h2c294c5890853e2b8400000000,
103'h0277be3a32989ee04eef8e8c80,
103'h16f245795ec1eb38e000000000,
103'h1c90b2fba039a9731200000000,
103'h2b51e8eaf92beeec7200000000,
103'h0a985d05d4bca1e81200261741,
103'h1e777000fe0e8ad30a00000000,
103'h11186e350aa6e7d8de38c32e16,
103'h22f315dc291e57d9de00000000,
103'h2ef9ac6fb936c60ee800000000,
103'h0cbce4eb5b29dbeb10defff5ad,
103'h2a8ea83a0923885ac800000000,
103'h1307536196e06d462200000000,
103'h229e5663016f15802c00000000,
103'h2b6c1f73557668e1c200000000,
103'h0e63c46eb614bf44c200422241,
103'h3b7ef1c4e280deb81600000000,
103'h3d7a8c6130e4a326ce00000000,
103'h3ee53c7dab6394ebb000000000,
103'h16c6557be6de214ce000000000,
103'h24bc2dbee4c35dca8a00000000,
103'h1432e4b9fa89b3467000000000,
103'h348e3edbde45e1055400000000,
103'h3e4d2de97378c5bf5000000000,
103'h2eea3e43e607049b2e00000000,
103'h024aac68e5543284a268e40000,
103'h1234cdd4523e70c88800000000,
103'h0364d04516891d316e45800000,
103'h240d987528bdeb05c000000000,
103'h2cbd65406a22bb4ad600000000,
103'h1ac164904f3053c00060b24827,
103'h1d03d4a8bcedb9006a00000000,
103'h32cf61f296af1d90bb00000000,
103'h3258da4232b2f2397700000000,
103'h1f050ddca682542c0c00000000,
103'h18e1953718db2e6e4000000000,
103'h0eabd591f6e03c4ae6500a0073,
103'h1a25337d8ec1d181fe00000000,
103'h1a5183a29d6da713f600000005,
103'h010027f3b892da9184c981429e,
103'h0089fab312e45e3422b72c739a,
103'h36f409bd54e48627da00000000,
103'h3b1fea49946e80daec00000000,
103'h1cb971e9ca628a984000000000,
103'h36e5d41b848274e1d400000000,
103'h24f69481623be6cb9e00000000,
103'h24ebdb0f1921bae72400000000,
103'h3a4fa277bd184f688700000000,
103'h1915f478a2042a779e00000000,
103'h3d5ebb5b5d53ccef5c00000000,
103'h02e36909b569c167fe00000000,
103'h2289d19f32c87cc35a00000000,
103'h3e48899d34abe5cd0e00000000,
103'h3c0b6c12d635b76c4100000000,
103'h16221b77d57e41097600000000,
103'h24a28c44d089ad1c4c00000000,
103'h26eb79d526abc8942200000000,
103'h1ce04d328c4e54d8f200000000,
103'h290ad7fc3339ceae1a00000000,
103'h0ab3a3cf4f1a1be0a600000b3a,
103'h3ee61cbeb724f3dcd800000000,
103'h18c45e4242d897ac2600000000,
103'h3ef0f49ec0beb46add00000000,
103'h175759a9588312ad1e00000000,
103'h3cd7da949674074bde00000000,
103'h197d4f5caccb60f53600000000,
103'h38fb5bd0e8a33b89cc00000000,
103'h16381cb000208ae67800000000,
103'h0ef7f03c381be6b76009f01a10,
103'h1b2bcb145154036762ffffcaf2,
103'h152b06e19e4bf3a39a00000000,
103'h34cd7e38b877beb7ea00000000,
103'h169080764ca2c5998800000000,
103'h336f696b437043d24300000000,
103'h1ca255c79800c4488e00000000,
103'h262135c78a702db3d000000000,
103'h2917d47f6912837b6a00000000,
103'h36b138d0ce33b942f400000000,
103'h08bae0f4764b8dc25c78b69b15,
103'h32c54d60acfcc6932b00000000,
103'h263fe780b4b7a787a000000000,
103'h04cd051c277cf4e84e00000000,
103'h2e8ddbfa8ebcdc690200000000,
103'h109a409b5289e1852a082f8b14,
103'h1ea36bcf4117bd7fb800000000,
103'h20643e8ad0b1fe1b0a00000000,
103'h0aa2062eae5569ea4a028818ba,
103'h029caa3b90b9a8751c47720000,
103'h0c212fcd9a5baea3ca3dd7f7ed,
103'h18bd72df5ef858df5a00000000,
103'h340bb40c2b1988acf600000000,
103'h3eaf5f2342d6fb8c5400000000,
103'h1a0cb2af76e2af987e00000000,
103'h10c5b4df76920ebbc219d311da,
103'h25770feed09ec16b3800000000,
103'h2341f3ab2064764aae00000000,
103'h24e3d2f3c4db86397e00000000,
103'h1e6861d4e61d79e49e00000000,
103'h0d7eff71cc014cd862bffffcf7,
103'h0d345e79eb69aead4abeff7ef5,
103'h2a4e33ccb6e8ae1f1600000000,
103'h0e438f59031d0c990000860c80,
103'h195664c9ee6b4065b600000000,
103'h2f6a87133caecfbeba00000000,
103'h2ee85809d5053488a800000000,
103'h254ed71f836fbb9be400000000,
103'h1ed262ce315813a5b800000000,
103'h06c12ee294a6eac53a00000000,
103'h2b5ecab5b5794d936a00000000,
103'h22019b117a3a7c75fe00000000,
103'h1d1427092699472bb200000000,
103'h067ec6a6889ae23d2e00000001,
103'h0690510926af09465400000001,
103'h381b28ff2c2dcfecdd00000000,
103'h26e07d6b32be20f60200000000,
103'h3b3f1902ecd949f53000000000,
103'h183896d7d2b9c7606200000000,
103'h1ae11df30ef8e0634e00e11df3,
103'h0ab774fb2731773b2200002ddd,
103'h2e4becf94112952e3000000000,
103'h3cb9aeec8cca0a295700000000,
103'h1ee138403a15f7229600000000,
103'h0e01a1f736cfa60f2200d00391,
103'h255382e956b0de4f5c00000000,
103'h3cb7f909a4b280469400000000,
103'h1ee679534b06032fea00000000,
103'h3d2af0bf86bdfc398e00000000,
103'h103f0e3ae4a4758cd8cd4c5706,
103'h3a040a05a0cf664c5e00000000,
103'h087b8616f10e748744baf948da,
103'h22f905582a127e8ce400000000,
103'h013480d2f48e04a3d6e142bb65,
103'h051471da968709fc0000000001,
103'h2ac3c92e96bb8acef400000000,
103'h00819509dccffca98aa8c8d9b3,
103'h0151df720693c5d822f2d2a514,
103'h36b02e7e07155ae1fe00000000,
103'h0095878607673a5404fe60ed05,
103'h22366b5cfd1768d20a00000000,
103'h20a74bdd7eacf0581000000000,
103'h24abf23620e35bb50e00000000,
103'h2ec5f370c28aa7928c00000000,
103'h00472eff663699c8ac3ee46409,
103'h0edfd36016fc8d396e6e409003,
103'h1b256818d743bc38d6fff25681,
103'h074e5886a5238f98ec00000000,
103'h3701f086ff48f7b1c200000000,
103'h0cec225004975038667fb93c33,
103'h38d2e1527a9940bf6400000000,
103'h3afd5c8dc685630f6900000000,
103'h204b6761ff584461e400000000,
103'h04e269e7f855a0efaa00000000,
103'h2c10bca658a10851aa00000000,
103'h10d850241c837239a22a6ef53d,
103'h3d2546b14a942edffc00000000,
103'h26ca81a05a6c7f041800000000,
103'h08c55d7f1691c5b5622a4c653a,
103'h046141af7d5c4755be00000000,
103'h1e8098198621a4d4d400000000,
103'h00341d638a82e684525b81f3ee,
103'h3e5421b1a9037e9dd800000000,
103'h1505ebb52a379c016200000000,
103'h2613fd0e688bbdb30c00000000,
103'h3e43b33c7c91a9683600000000,
103'h20f64feee2a5a6769e00000000,
103'h2cac6b3f20e959b31c00000000,
103'h229a2290c2dfa9a1fe00000000,
103'h021397956e8c14e120cab70000,
103'h1f1eb60253263771e200000000,
103'h1ccf7ae5d439cf075000000000,
103'h3d69997c72588509a200000000,
103'h1ee361b50e27ffef7600000000,
103'h30e93ececc91996be800000000,
103'h1215535a6b74fb20f800000000,
103'h0a7b36ed5b5e39efc40f66ddab,
103'h33399f89ee738d4a2f00000000,
103'h2b200815f8eec4378a00000000,
103'h2e980a0deb2863c17800000000,
103'h1e850726d7486bd77000000000,
103'h28d03e2f84e075e55a00000000,
103'h208f028262657d0c3000000000,
103'h103c8b0ccb35bb3bb68367e88a,
103'h2a127758aac4bdbe1800000000,
103'h1c30cf7bfb0148cae400000000,
103'h132f9d84a613c0238e00000000,
103'h2a93e89983448f9f8a00000000,
103'h0f2deeea15742d243092161008,
103'h1e8cb2f8bf0815bdb200000000,
103'h28ecbfd24f3604a7c600000000,
103'h19608ccf6cc2b7a08400000000,
103'h0b18e96c14af7772d200463a5b,
103'h1145732cec1004423e9ab77557,
103'h157a12ab7628edae5200000000,
103'h28e4b6d1c66e60db3e00000000,
103'h261212989ae87386b400000000,
103'h3aeee5d242cd2a587b00000000,
103'h38dbbd4e2adf3cf11700000000,
103'h2ef1827864ce22c35800000000,
103'h2875a87ddca9e0118200000000,
103'h3ee2420a0a9b6289e700000000,
103'h191c05eeb5110b07c400000000,
103'h1a3506c472f34d11ce003506c4,
103'h021c2a5d8a0f5300821c2a5d8a,
103'h06ad2e08274459c4f600000001,
103'h14d9943ca86084228000000000,
103'h19170578ee0db22aa600000000,
103'h0e47c3c702e746674e23a12381,
103'h0e87d5159afe4be03c4320800c,
103'h360c402929460fa74000000000,
103'h04f12f5f38cde4bcda00000000,
103'h02e3d0bfeeda24e604c7a17fdc,
103'h02bdb887f2cb54453c40000000,
103'h1c95ec3034af25052a00000000,
103'h20b42f7fb66cdd8d1c00000000,
103'h1ca0578c1502c9bd5200000000,
103'h0666a47e74b6f93d0800000001,
103'h24f845b6125750c91c00000000,
103'h36390bf2d8bdf5479200000000,
103'h3ee6afbcbcb63afda500000000,
103'h1c971d43f2ef46f07c00000000,
103'h2efe840832d5f6ad3a00000000,
103'h12bd3b958e6d13f12c00000000,
103'h0f39e86a7c6b97f95e14c0342e,
103'h096cd03d0e28d38eeca201d9f1,
103'h368eff001c62bbf96800000000,
103'h1487247066cf8c367600000000,
103'h02ec5dd1dd5e8b3694bba3b800,
103'h2abd2f2cb0e5afa6fa00000000,
103'h22b6d41672d20d78d600000000,
103'h371334f99e8f3ca58600000000,
103'h313f2213414610bbfa00000000,
103'h06c99a63775945b59800000001,
103'h0d39c25aa69867c8d8dcf3ed7f,
103'h077bf7caad62022c4e00000000,
103'h1e4d69e0389bc486f400000000,
103'h3764ecb1c117bc51a000000000,
103'h04d5b538de652631d800000000,
103'h38dee588d6ca12e39800000000,
103'h184a18051a9fc81c7800000000,
103'h33510f08557eada54f00000000,
103'h0a6fc25d2cc8c5aa680000037e,
103'h02f39be3de19d4b2bcc0000000,
103'h1141884e2a89970fea5bf89f20,
103'h3a2f3cd4ec7d32f3c800000000,
103'h369b9f00febebb41f200000000,
103'h20d0c6d778edf816e000000000,
103'h2a1fc360ae899717de00000000,
103'h1cf856f9d15a5def5600000000,
103'h3d4e1d86ba7a21500400000000,
103'h1a629f5596727849d4000c53ea,
103'h3165193b54c095d08e00000000,
103'h36f12a38ef2335262600000000,
103'h0ad79925e0884e617a00000003,
103'h1b382962d679789a68fffff9c1,
103'h000b31e9a05111c0482e21d4f4,
103'h3a9ed040fa893b231f00000000,
103'h2255a3be7a946d0cc000000000,
103'h2c94c59d74333d4dba00000000,
103'h0b4d6016d888e10c3600000014,
103'h0b570c50841da6a9aa0000055c,
103'h06e9f3ad4e6b06c08200000000,
103'h3d114816dac213110600000000,
103'h276bd9ce20ac06be5600000000,
103'h2b4f4c919cbd4ed53000000000,
103'h305065fec32928a35000000000,
103'h06bc862c6d787534ec00000001,
103'h36eab96b1ec8db33ae00000000,
103'h06c4f368248561601c00000000,
103'h335c7c3a5d701acb3b00000000,
103'h221d2dafe2350e335e00000000,
103'h3f56545a56918a6dbb00000000,
103'h3958563878aeb81d9f00000000,
103'h16dfb976b7050c77f400000000,
103'h12d737802f5d62b06c00000000,
103'h3003c3bd053d1c272200000000,
103'h24c1da67971453a75000000000,
103'h102ea92fc6181764540b48e5b9,
103'h32a0846fead9f1cbed00000000,
103'h026fc2607a089afbb27a000000,
103'h167c1c782ca91f6b9e00000000,
103'h029cca372e18e1cc1851b97000,
103'h36d58f5a8694fe444600000000,
103'h14e84649c831c87b7400000000,
103'h2c039834be0757d5fa00000000,
103'h32c8098b52ef9e1fc500000000,
103'h28a55cae00f336548200000000,
103'h2217ae14f2bb3fdfd600000000,
103'h26bbc7f75b609c8dd600000000,
103'h2b6739afbe784aa2c800000000,
103'h00024987e534129a249b2e1104,
103'h16908fb48e9b4c49e200000000,
103'h1eda15c10e9d95d1c600000000,
103'h0284385b652e258656e16d9000,
103'h24a6a59884083b476400000000,
103'h2cfd256fc68c73a2ca00000000,
103'h02eef190ed33193b4ebc643b00,
103'h277e5383d8303eab1400000000,
103'h313bdafd1a1f303c0000000000,
103'h3e019dbdc09d83bfd800000000,
103'h1553d42132d95ebcf200000000,
103'h14d923bff0dafc7ab400000000,
103'h2e8eb209c52ed09be600000000,
103'h2163708f9a07f45bd600000000,
103'h14d5b2d54896a6659c00000000,
103'h3a2153d7e8fa16f53600000000,
103'h1347f1553ecfc9ca7e00000000,
103'h2e9d5f6e78f11da26600000000,
103'h24fac1e38a390ef7a400000000,
103'h22eecabe38d66e661e00000000,
103'h08dcea8e1cd13049a806ed63da,
103'h2e9ad4287ebffb07e200000000,
103'h0d49db65489ce595feeefffaff,
103'h3531f199b737b9be7e00000000,
103'h16f0763442819523c600000000,
103'h16802b1876b386bd7c00000000,
103'h14cfdb048ea3fcf1be00000000,
103'h1abc7086a424280a3400000017,
103'h16e0bfc738f4030ec200000000,
103'h1486a42b92b073956600000000,
103'h08e00f4d6891335c9e389e08fb,
103'h0cdd7760fc17d788306ffbf47e,
103'h32ff077ec4f7e6d59900000000,
103'h12149aab50d55e369400000000,
103'h02daa16d44d465b55a16d44000,
103'h1d31db8bd6e90060aa00000000,
103'h30a0ed3298c3a1cdee00000000,
103'h0a07e5aef4f57d59c400fcb5de,
103'h37443c61e6966a8c5e00000000,
103'h2454f8ca309e503b5200000000,
103'h2a4eb59326e28c9d3800000000,
103'h090c142a0d3785676a1dc8a6b3,
103'h1abef01ab6863afa90005f780d,
103'h15083697be924f249c00000000,
103'h3eefcd5018513f3f5300000000,
103'h0eb9f0a5ac5975d7100cb84280,
103'h2cbb9962ab4943272a00000000,
103'h3f437d1a3a0333ccd700000000,
103'h115daff666becd2f824f716372,
103'h3ac92211e5024a49bd00000000,
103'h108e0a04755ffa40229707e229,
103'h129c351e2e291c520600000000,
103'h0ead9404c0b726567c52820220,
103'h307dc01ad2535b74aa00000000,
103'h3950367aa200ef796b00000000,
103'h3482a71a937eaf943e00000000,
103'h1ede340c8acee60ee000000000,
103'h0af0e754fe518d29720000003c,
103'h0956f6121f2fc135fe3c9b93f0,
103'h28bdf448a820a88afc00000000,
103'h1aa3a21370779e9d1a00028e88,
103'h195835ed183592e5c200000000,
103'h165e56f032d934f93200000000,
103'h309439294c316ae64a00000000,
103'h34eac3ed628fc1d67e00000000,
103'h26b8ed4e9323faffca00000000,
103'h32bca995870ebeed2d00000000,
103'h30999ad5aec7ac3bbe00000000,
103'h3aa7f6fc208455d14700000000,
103'h274614f9111df0a6f400000000,
103'h25082df5cac5e7a31400000000,
103'h2ad905dfb10bfc9c2400000000,
103'h1e718a0555142a91ee00000000,
103'h328e63fc40ed30719f00000000,
103'h16c92e9a1e5eba76f200000000,
103'h04c9e0db12ed1e733200000001,
103'h22d68fb828b64d0d5200000000,
103'h16f769272e802de86400000000,
103'h08057307d056bda08c29e753ae,
103'h1a72375f664e26c7ba00000001,
103'h3ecc1a2a315399cf8c00000000,
103'h0cdc4a024ac5d12ef26eed977d,
103'h076ca7c2ca91eb592200000000,
103'h1353c323d76e355b6e00000000,
103'h0689054c9cdadd1e3800000001,
103'h2911e144f12ea0420e00000000,
103'h17608e6c36b7a58eaa00000000,
103'h0e4126ec9ec986d39a2083604d,
103'h1c8ff4c8762a153fd000000000,
103'h08b99fc2856b3c2c70e951f77a,
103'h2311eafea2fb30f4e600000000,
103'h3521dbc96ab4d0b76a00000000,
103'h24fb5367ccc6bbb60c00000000,
103'h0afee04600e8977f760000000f,
103'h346da950a4e3eae74400000000,
103'h02d7a3502ee2cb2d44af46a05c,
103'h38f66e072550747dea00000000,
103'h3cdbf474262817ce1800000000,
103'h02aa12609e1e85d53cc0000000,
103'h2d5c1b345cfa7a496200000000,
103'h04f0ef355ea48caa0200000000,
103'h02d637b44b00a7de5eed128000,
103'h24e398014ef19713bc00000000,
103'h260f7e2390c7cec80600000000,
103'h0535de8f36ab66c95400000001,
103'h0000cba4dcbae4ece65dd848e1,
103'h06cc6098e2f0c37c1c00000001,
103'h1c898ca0a2f18f20f800000000,
103'h030e87706abdefb9da7706a000,
103'h1f3ee90987477c5a7e00000000,
103'h172a2f8f895603cae800000000,
103'h33063991a694ecd46f00000000,
103'h30d3d2b4bcbf1c63f600000000,
103'h185f5b91aec555f59c00000000,
103'h063260c91e9928aa5800000001,
103'h3c5b69cb76f8843c0900000000,
103'h18195fa23c2ae5052600000000,
103'h309671dcf8864ed09e00000000,
103'h38d8da0d509fae72da00000000,
103'h20b46ae80336204fd400000000,
103'h3e887ffeba0efa5d2500000000,
103'h18877a1a9ac365452600000000,
103'h2c0cc307194be543e200000000,
103'h1331ba6672d35f5e7c00000000,
103'h388cd2159ee022659700000000,
103'h1af6e421f111dccc0807b7210f,
103'h19245b736a9eaee1a600000000,
103'h2e9db808c49593039800000000,
103'h36ea73fc9cb9ee770200000000,
103'h1c1752560a57a67fc600000000,
103'h34560d7b81421a7c6400000000,
103'h373377829e596cd26e00000000,
103'h3ea6748d52af7a4df000000000,
103'h22d3600f0ae2f1d08e00000000,
103'h1157f2108889665de06745d954,
103'h011e9e8e6a5cc66ceabdb27daa,
103'h0e3eb7debab4b87d721a582e19,
103'h310e4b7cfcd3570bdc00000000,
103'h1ac0d0ebcb120eea9800060687,
103'h0efcbcb87b205a6794100c1008,
103'h2a956ef216e12b535e00000000,
103'h02e2d9a924dde80bda9a924000,
103'h16039b6c0f7356fdf000000000,
103'h37366c19935630a71400000000,
103'h1089972ea859cc132217e58dc3,
103'h00bded971e90382cb4a712e1e9,
103'h14d02c0b6f19cf5b5e00000000,
103'h3655c17daed7bcf27c00000000,
103'h2c31879702a7e8fdec00000000,
103'h0b6719c37afdaa7b9a00059c67,
103'h072ce41ca72f32129e00000001,
103'h330c7dd130964bd61900000000,
103'h0ec3d47836c32ff2be6182381b,
103'h2d23141d2acfadc3ee00000000,
103'h057ffe3db893823c2400000001,
103'h030c1a70e4b696594e069c3900,
103'h312e827a283694970600000000,
103'h15141a762a42af07ea00000000,
103'h24c960361a7131821200000000,
103'h2a1228322e854bf83c00000000,
103'h16118687924eac2e5600000000,
103'h29477973ff60d4608600000000,
103'h26c01b6854725ae81800000000,
103'h3ca9eedebcb9d45c1700000000,
103'h02190e4d6279efc46ad6200000,
103'h1cd6d9ea6123dea32800000000,
103'h32f579e7e23cecf08b00000000,
103'h1e8674cd7e13c6daea00000000,
103'h06d1440f330940c2ce00000001,
103'h10960315508fb5904c0326c282,
103'h3d7ea0be9660f99f7e00000000,
103'h0aa42b5866f6fcb4ce00a42b58,
103'h16dd7ccd22759d736400000000,
103'h16200f04ad19c8cbcc00000000,
103'h24f256cc84f74598ee00000000,
103'h0b259833db17549d9c00024b30,
103'h164fd64fff09ab6a2000000000,
103'h04efb1df892f439dfa00000000,
103'h20a9563ade7f19edf800000000,
103'h015a402f256ecbcd826485fe53,
103'h3a227ec1041822086100000000,
103'h34f468bd067262378400000000,
103'h36f596570094e0f88a00000000,
103'h1675dddef48949b59000000000,
103'h1c64f1346a7ee00c9000000000,
103'h276c269242f4bdeb8600000000,
103'h36e5be279e59af1ff000000000,
103'h06f436b584c5d5b23200000000,
103'h0c8bf8f8faab93d9d055fdfcfd,
103'h3ea29b49009fca8f5500000000,
103'h30adfb848e2bc3884e00000000,
103'h03130ae00cce5ed15085700600,
103'h163defedbd7c5a55de00000000,
103'h261468d53e8f6535ea00000000,
103'h368aac4c16cd5523a600000000,
103'h152cb34b3ce1bdf8e600000000,
103'h3e9d191bb36c6a44fc00000000,
103'h2489d94206991d903800000000,
103'h0b05fe9e453636abea00000417,
103'h064f791e28c00fedf000000001,
103'h3f7ab196f4c60e8c3500000000,
103'h28125454ba1587aa5c00000000,
103'h194314a2ba9039415000000000,
103'h0caa0b9ca2a28d960c5547cf57,
103'h2ad112847ce5a238c600000000,
103'h3abe27f8888fadd56900000000,
103'h06c0c516f260c059e400000000,
103'h0d539b76af1ee8526eaffdbb77,
103'h3688ff6c74dfad696000000000,
103'h1aa4059b023348e00e00a4059b,
103'h094eb99ef8bc484c84f978e93e,
103'h2a5a2dfcd3604de78600000000,
103'h38848aad1caf07867f00000000,
103'h3c8e94c6c60935835000000000,
103'h02cbe7c07e8dc0306c0fc00000,
103'h00c58306bc1c54f73270ebfef7,
103'h121f6c347ee83cb7b200000000,
103'h3f285ce8c0adbfbe6f00000000,
103'h333a832052cd2bf2ed00000000,
103'h24da698850f588dbac00000000,
103'h1296a4e782300bfbfe00000000,
103'h3e3b1cfe670a75845000000000,
103'h2c8d54d3b8a11a6bd200000000,
103'h2aacb89bf8dc376a3a00000000,
103'h3ac1a53fe4698c3df300000000,
103'h0e069ddfce1644d9ea03026ce5,
103'h09560c040ad7ea19cec0f30ee2,
103'h3b46949418de87f99e00000000,
103'h2713548e613493fda800000000,
103'h3449a0c69b7b2891c000000000,
103'h129631d8c08e7d202000000000,
103'h3abaad04b6d81de6ba00000000,
103'h3abdb02a496e4fbf7d00000000,
103'h1af5474d8528fcc4320000003d,
103'h16a807027ee6acee7a00000000,
103'h12e943d79adbf43bfe00000000,
103'h05029e937083fb3e7e00000001,
103'h3e8a490ec36d3f161800000000,
103'h3f3af04e476fdda98800000000,
103'h3cd2447c44fa26b84b00000000,
103'h14458ce6433517069000000000,
103'h1c3cd08ebe075b82d400000000,
103'h26a1534d534ce8691800000000,
103'h3675b3b56e89b8f7d600000000,
103'h0a443ad5d52b0c452a00000110,
103'h2247d8fccaa0bffa9800000000,
103'h3b52d2a696e4fad06e00000000,
103'h24aab4b9782cd3cd3800000000,
103'h3c8c4fc4327fa673ce00000000,
103'h2a98f714172a5b2d4800000000,
103'h25465e5e94b6aaf17a00000000,
103'h32d8c0797f4fa2059300000000,
103'h3a97f661a29600642700000000,
103'h36d6d2bd966ec0dda400000000,
103'h08400a46d106b73f48a35ebccc,
103'h2e5fecc186dd89fcde00000000,
103'h12cf7141ce1d9443ae00000000,
103'h1ad4f6263d7d8105360000000d,
103'h39493be8504cf2470500000000,
103'h28c438e9ab21e86d4200000000,
103'h1f1cbfe7e56b24559200000000,
103'h2292db29cc2f5d3f3c00000000,
103'h24867770ea4c1d272000000000,
103'h36c705ff0cdef850ec00000000,
103'h35297cfa72656fc1d600000000,
103'h14f7184b692c75c0e400000000,
103'h02f410db9d55f2bb56436e7000,
103'h193d2692f24d0b06be00000000,
103'h3d65349b35411be25c00000000,
103'h12f2b2654d7e42754e00000000,
103'h12aca5f04ae377108200000000,
103'h2ebc8c369cd62975ce00000000,
103'h3c197d83ae82cf661900000000,
103'h3eb78ab31d3f5b9cb600000000,
103'h0cd3da57d858d920646dedbbfe,
103'h26d3a10d171063d38200000000,
103'h1ca9913824e43e2b5a00000000,
103'h010250c94ab7df3872dd1800de,
103'h029a6bf72761707096afdc9800,
103'h1e8b60456763c139e000000000,
103'h108cb8672afe2d3106c7459b12,
103'h27724eb448898d766c00000000,
103'h070fc439d81645dd9600000000,
103'h0d0eaa2ffe889491dec75f5fff,
103'h39715160049858cbb700000000,
103'h10d225c110a702fbb4159162ae,
103'h2ebc87988818545bb800000000,
103'h26bd2f4d98ea7a1cc800000000,
103'h1b466b9488a701b552ffd19ae5,
103'h156800a72e643102ea00000000,
103'h1c3098b588aa9c977200000000,
103'h2e11851f9c129d3ea000000000,
103'h1adceba67b4335f42a00000373,
103'h0c4f53e2a854bb13c62ffdf9f7,
103'h2e25ed21c231a6ba4000000000,
103'h18a722f85080fa9cea00000000,
103'h1f3af60d7ea6e7beac00000000,
103'h2111ff16d64e0ab6fc00000000,
103'h0a3dc333f48900c47a00000000,
103'h369b2e0b549affdb5000000000,
103'h3479937f9ed8c30f4600000000,
103'h2efee0b29673f11a9a00000000,
103'h00d2389c8aed849a3adfde9b62,
103'h062e914af8ec654cd000000001,
103'h2025e9d4b8be9de95a00000000,
103'h1af6056dbeed2f3452003d815b,
103'h2b3a1221611319090c00000000,
103'h046ba36f3a091e76ca00000000,
103'h18899a09e64330982a00000000,
103'h24662e8deaaed4076600000000,
103'h2e2ff24643386e114c00000000,
103'h1a0ccf07a69e9c9f3600000000,
103'h00f2ca3fd6ce8ee57ae0ac92a8,
103'h0d1bf61030db5ded20edfffe98,
103'h02f3f5e7f0ce282cf6c0000000,
103'h3d0463d0fcea1e3d2600000000,
103'h1eb36e593ede14251600000000,
103'h153107c6fce277f61200000000,
103'h3c89ff21da95e64f5300000000,
103'h12b11ea9aec6ee164e00000000,
103'h26c25c6eab50ed382800000000,
103'h38b1ae58be020be1d600000000,
103'h06837838e4c468508200000001,
103'h2eeb28685d7616a94000000000,
103'h0519c6ae22f98ee22400000001,
103'h0699522c10e4b74a8000000001,
103'h061ae98bd4fe7df8a200000001,
103'h2b60e93c1c97d024b200000000,
103'h2a1cff95a2b2b9b08600000000,
103'h0cd2a4d14e13a2eca269d37ef7,
103'h3e6d01577930a2824600000000,
103'h0705dbd6470347539400000000,
103'h28368679c47048ab0c00000000,
103'h2e19eacdca7624815200000000,
103'h0310f20e74acaafb189073a000,
103'h10389bd162c695c8e2b9030440,
103'h23638ce7e6d787d75600000000,
103'h3afec6a9771023a8bb00000000,
103'h1e1024ec5973b090a000000000,
103'h34ce2e2a5572773a1600000000,
103'h2f52cd3132829c266e00000000,
103'h0eaef40f6650ca50c200600021,
103'h251b3e9656a39781f400000000,
103'h14fb39ade5528b915c00000000,
103'h174dabff8b6dca27b200000000,
103'h0d22ba779e6903d596b5ddfbcf,
103'h2848934074b6afd52000000000,
103'h1a12038b40d96a4cbe00000000,
103'h302dff676921fd8d3400000000,
103'h12b7c56b423401187400000000,
103'h10aa8f44b562007fdea447626b,
103'h055408f34619c5eb2000000001,
103'h3ad6ecee96c4552fd500000000,
103'h197bce771c185e231a00000000,
103'h3954b11816ef4b11b300000000,
103'h0e8f9438ef6b1988ce05880467,
103'h28e43d44e6bfcaa0e400000000,
103'h1afd3b80b54f5ed9d2003f4ee0,
103'h292e97df9e339c1eb800000000,
103'h0c4f3f503930d79f6ebfffefbf,
103'h1edb0049a35f6f7f0c00000000,
103'h18268be3eeaeaecf4400000000,
103'h06c176580e89af18e600000000,
103'h128ffceae6b03afcd600000000,
103'h168f5b1d2d71b154e400000000,
103'h3eee28ce7f01ae3fca00000000,
103'h14fba54f1491095cf600000000,
103'h3892d0e8937f322b7400000000,
103'h02da377ee67ad77a88d1bbf730,
103'h38934f6a1f0da8631c00000000,
103'h2c4e159520e7dfe20200000000,
103'h3499e51d197b2f4c2200000000,
103'h1064e6d084c944e142cdd0f7a1,
103'h14aabffe7b6329fe5c00000000,
103'h36fe418f8ac810cee000000000,
103'h3839a3029e72d0cd5b00000000,
103'h14f033c1d571125ce600000000,
103'h377009624eaab55f8400000000,
103'h10530901229ae9215adc0fefe4,
103'h36fe196ed90af283a800000000,
103'h3d1bfaa9ea5dfb84ca00000000,
103'h16aaee41e15c14f3a400000000,
103'h3ee497395d780f9d8e00000000,
103'h08b929523222fddf6e4dea46ae,
103'h2c98adeeb1079518cc00000000,
103'h3ad62e0ffac0be6aff00000000,
103'h2a6fc324e7596c59b000000000,
103'h368167d7632f9a69aa00000000,
103'h34b60a694c9f5d8e9000000000,
103'h24f242140220c565f200000000,
103'h0eef3829b6d6cfcf3e6304049b,
103'h21459a991cc911e34000000000,
103'h12cb97722ab84a0cf800000000,
103'h12f0f1d9cafde4a61400000000,
103'h133711a75ec97c183e00000000,
103'h0b54014430ba6df20a05500510,
103'h1e3a02c442f17f996800000000,
103'h1ed84e514f4580dd9800000000,
103'h28747e846c7f83a1da00000000,
103'h10da2acfca57d1f328412c6e51,
103'h28fa450d32cc50779600000000,
103'h020bdee402a67b476072010000,
103'h2c62f9986aa0c0549400000000,
103'h033997eeaeac9f38965fbab800,
103'h236808381b0f98d10200000000,
103'h3762c8f91d4930bfb000000000,
103'h0e0405017eb138f7ca000000a5,
103'h1146015e771401f0e618ffb6c8,
103'h01349cf4041806f264a651f334,
103'h0b32d15a945e0850da0004cb45,
103'h317a3680d492a544de00000000,
103'h1572d49edec5769f7200000000,
103'h317f74adce3fad204600000000,
103'h0ea41baf22b281bf245000d790,
103'h0226cb015231f66cf252000000,
103'h093c1f9862d6121c16f506c23a,
103'h2f16eacee4fcdd1d6800000000,
103'h20316325ac38fcb5ca00000000,
103'h36fe5d3b9a4fe784ae00000000,
103'h20fd4dbe7c814aaa5c00000000,
103'h2ad2505d727fa7e5f600000000,
103'h1aa43019d27cf5a47200000029,
103'h36af0c8bff4f4601e600000000,
103'h2d09d082d8f3761bb800000000,
103'h20e5df240ea282a7b600000000,
103'h064195ab3aac532a8e00000001,
103'h3e1a41d6da92324e9c00000000,
103'h3642340460d3c7f9d800000000,
103'h055d9c4da0ee09d0b200000001,
103'h231b873e97303dd51400000000,
103'h3a85c55a1a8dda22b400000000,
103'h2c8235c43ca961614a00000000,
103'h00526e28362f26bb6440ca71cd,
103'h3510b05ce4b15c7fa200000000,
103'h3eff3066a403caa7d900000000,
103'h257b8a931a147b04bc00000000,
103'h06a14620d913ab6b6200000001,
103'h1ef62869fc8f35fe7c00000000,
103'h1cfc6732c2307c1f5400000000,
103'h3f0670a36326a4895200000000,
103'h3b24f518be230bbc1400000000,
103'h0f5724f97c297c5f7600922cba,
103'h21188ad8b64e71783400000000,
103'h360a6cd744a59671b000000000,
103'h2d22f35f26be214a6600000000,
103'h235e85a31cc88e21ac00000000,
103'h12c3944688eb8180d200000000,
103'h3a7714622b4a0723ef00000000,
103'h26d02aef7e0d9b6a7600000000,
103'h38e762c73884afcca200000000,
103'h26c728c09f54dabc2000000000,
103'h1c92703ad73c3d835800000000,
103'h3ea7bed8fd036643f600000000,
103'h1ecaa8e19895d67ecc00000000,
103'h377242b6d93d9557c800000000,
103'h2c6eb74836083e396000000000,
103'h38a7695cee7a80f03800000000,
103'h00e381b59ae9383870e65cf705,
103'h22b5708d1490a1955e00000000,
103'h1ac4f4bc5474234af800000006,
103'h0adcb724f62993d80c01b96e49,
103'h296efa7dd2ee88946200000000,
103'h22ea760f1ccb3fb95800000000,
103'h2ef69335c63a3a372a00000000,
103'h1176d3a76924b046482911b090,
103'h2a20a7f1171b437c0e00000000,
103'h14b904cf289217237600000000,
103'h1d1ca16692b2bf148c00000000,
103'h2aba7835266bc3e3b400000000,
103'h217cff4a0488654a4600000000,
103'h2e5ac9daef42dd7f6e00000000,
103'h22caab8f50bfdcc97200000000,
103'h2aed4c583e1aa6a46000000000,
103'h187bb104e0e55233b000000000,
103'h0a927afbcad29e8bee00000092,
103'h2aec2272234e4f90d000000000,
103'h1c05a6b1ece0ca8c9a00000000,
103'h0b39d19618ccecfebe00000001,
103'h1b534eadf4d293b0aafffffd4d,
103'h363f6a51be0c6546c200000000,
103'h3579d5865a5fb3f4b600000000,
103'h1e950b47909f1e467600000000,
103'h237d2e078518f3ccd000000000,
103'h1837e47822adff146000000000,
103'h0eff002f852b2d1be4158005c2,
103'h1f25cfdb9e6311940600000000,
103'h3eebbdce2d6211c38c00000000,
103'h22ca9f8d8c87e19f2a00000000,
103'h2a5780614a739f6d5600000000,
103'h370f8e50ee3e3efae200000000,
103'h212aadd49895bf5c2e00000000,
103'h36a7df1bcea54dad1c00000000,
103'h1aacf2022ecffb81b400000015,
103'h0825a455e577da9d82a93f6433,
103'h24dc95a47f24cc9fb000000000,
103'h1829464f464a70f59400000000,
103'h1a1b44a72b27069a1400036894,
103'h0add3e80c2504ce95a000374fa,
103'h1e1712f7dd6b91908600000000,
103'h3275b40ea648d0114900000000,
103'h0f1ec61b075fe309268f610483,
103'h14eedec178d59717cc00000000,
103'h1c0f445146f45d32d200000000,
103'h029b3b719ae33bf44c676e3340,
103'h117002a338f28045923ec12ed3,
103'h22a4acddfa8dbbb72e00000000,
103'h2eaeee308afdbe5a6600000000,
103'h02ad8cb5eea26b38605af70000,
103'h308f672f9d515968ec00000000,
103'h1663c1eedefee61eda00000000,
103'h36c5d8654e8e4d4e7600000000,
103'h2225ad3624f20f3d5600000000,
103'h3d27ed3f5cb7e7a2a400000000,
103'h347b86b17edd94d8ca00000000,
103'h0ace06427d0582182600000ce0,
103'h2eaed321f08108c9a400000000,
103'h3881af3eba4f0f0c2000000000,
103'h1e0c72fe28fde22e1000000000,
103'h0574cb96627f916cca00000001,
103'h24e2a646c08c046af400000000,
103'h36d189c0c500d0015600000000,
103'h010f7c46eae3764816f9794780,
103'h354b50fb20b50008dc00000000,
103'h0a06b71c20c47c4fc6006b71c2,
103'h234e21a8170fcd4ae600000000,
103'h3e965c35601684670700000000,
103'h04c20d0ac264a60f1c00000000,
103'h2aa2bde900fb02447e00000000,
103'h3047eb1704bd0f4f4000000000,
103'h0efce58fef5fcd38422e628421,
103'h0cc8646fe0a7b84f4677fe37f3,
103'h0cf8895eeea49ddf367e4eefff,
103'h0f23b0927b6d024f1690800109,
103'h160be71547658bae0400000000,
103'h0d53ead056893c407eedff683f,
103'h2343a6daac952355c400000000,
103'h26d800c438e90e261a00000000,
103'h24d95cfcda2cb500c600000000,
103'h294044e38004b5c4fe00000000,
103'h0530690aa4de12c1d800000001,
103'h0ab5b0878c1e57a5580005ad84,
103'h0a24062a904ec0affc00000000,
103'h22bf10ce5d0471378a00000000,
103'h3d5ed137262877621a00000000,
103'h38dca461c8e788307700000000,
103'h0278cf31c44659679ce6388000,
103'h1f63bab1bf22fdc96600000000,
103'h14531769409bccfb2a00000000,
103'h326aeb82deff87ace900000000,
103'h196a47ccf5529f162a00000000,
103'h02affd7ea6bd8a99087febf530,
103'h2d18b0f9be27d265fc00000000,
103'h161d317000d7cfe4a200000000,
103'h1e2139932cf080de6000000000,
103'h1c77e0cc830db24e6200000000,
103'h3e8c129ee22eebe18f00000000,
103'h20c816d73ea6ccae1200000000,
103'h02dbeaf43d32df4cf478000000,
103'h10e03fef9cfaf62432f2a4e5b5,
103'h22f247395ed6e1186e00000000,
103'h17333a64b0b721080c00000000,
103'h081afa3e12a968416a59c93fbc,
103'h393599646adca2a61b00000000,
103'h044b2eaef2f79ce42e00000001,
103'h2e37a511eb2d36489800000000,
103'h0adb3c7cee7864f78a036cf1f3,
103'h39283c295eb00a097700000000,
103'h1151de7be88b468664634bfac2,
103'h1b731db2a0b382afc2dcc76ca8,
103'h10c19331f005612baa5e190323,
103'h36886da8ca787ede4a00000000,
103'h38ff52291c3a12103a00000000,
103'h25017d2fd2c27fb90600000000,
103'h2eb72ae64ac1d1e22200000000,
103'h2a7239c86ec34f11f400000000,
103'h30a5c788de7a79f83e00000000,
103'h1313675988ecb3c0ae00000000,
103'h074386e338927b498c00000000,
103'h0535784f0aa5e2a31400000001,
103'h32eab8ccd0e969864d00000000,
103'h3e1a7342d51ee1d55600000000,
103'h1336e17989099aa22600000000,
103'h1ee5caf9c6240de4fa00000000,
103'h353a971d1a5aef5e8200000000,
103'h1a78ccc6b940ba584a01e3331a,
103'h16d5e445af7b51756400000000,
103'h183c9666c8f41e3c1c00000000,
103'h22c7566cdeca0281ca00000000,
103'h06ad05d1790698e89400000001,
103'h24d36f8e5acdef557200000000,
103'h2f752ac0a27af526ea00000000,
103'h030b042f074e64b5462c10bc18,
103'h366ae01f34c38f75e800000000,
103'h20d154f7f8ce93a4ee00000000,
103'h2705b9262e3973c42200000000,
103'h0eb5127b4e0ac8bc1a00001c05,
103'h3cb2d085b61081e24800000000,
103'h20741e0604c5945d9800000000,
103'h3b03ff2b437864e34e00000000,
103'h04cd5414a2ec82e95200000001,
103'h1ca171ba1cf082149400000000,
103'h2a861141e0bdd6293600000000,
103'h3c3045273d5f47e35500000000,
103'h1252ddefe6e559253400000000,
103'h0961f9a1e5159e4c723a33f6cb,
103'h1d61976876687c3c5800000000,
103'h121f0b583eca75de3c00000000,
103'h053bc72b5c2c0d46b200000001,
103'h1d3ddc23af4b189ef200000000,
103'h1b558f687286dfca4eff558f68,
103'h0cd5bee98ec4bbedfc6adff6ff,
103'h3e206448e91a4b566e00000000,
103'h0c9716eef6f00a3ffc7b8f7fff,
103'h0858e233f5106e88e6a4465d89,
103'h36a18d4342a78577dc00000000,
103'h34aef4408a0067abd000000000,
103'h1ad6a69442a1f4ef120035a9a5,
103'h36ee6327f750e92f9e00000000,
103'h07168e4491278fc3e000000001,
103'h1ae63ed90715f2ebd6000e63ed,
103'h38b657194d2c81306600000000,
103'h18286448a712c0096c00000000,
103'h2eeb5aa79ec91722b800000000,
103'h14d5e0ca76f17b6b6000000000,
103'h00d659d924dcd612fed997f611,
103'h3803541838b2b6dd7700000000,
103'h18430e60b88910b69a00000000,
103'h194bdfcbf28c64ced400000000,
103'h0e462ca28acf732f8c23101144,
103'h281d4f8c221b52fb7e00000000,
103'h3ca7295331617f9e0b00000000,
103'h0aba13d0da7ecf2a2c00000174,
103'h0859631d5725f87d5ebe4db004,
103'h12c8259960e00c4e3800000000,
103'h01523b10ea396f6b8ec5d53e3c,
103'h1e3dd0267d019504f000000000,
103'h16a834663d53d015da00000000,
103'h243891235a91a03c5600000000,
103'h14a8fa2eb139d4a29400000000,
103'h2f52d2a5967265c5ee00000000,
103'h06fe40216b1b5ff4a000000001,
103'h1afd7db31b6e329a360000000f,
103'h088e5b81206c72bba071149d40,
103'h29590df1ba69f06eba00000000,
103'h1e96262842f84befda00000000,
103'h00ee9e536c5159e1949ffc1a80,
103'h3ab54918cae78009d800000000,
103'h16e86699cad61e5d4400000000,
103'h2a857489868b67760e00000000,
103'h031ace691d73ce0fdae691c000,
103'h0601822a46f942996000000001,
103'h16cfb5f54b1411027c00000000,
103'h3074081d9015932cc200000000,
103'h10a3c1bbe6e549220cdf3c4ced,
103'h0c47496a1759513f9eafacbfcf,
103'h0ee413b1a6fd12fb84720958c2,
103'h1c94eefbb3445c659c00000000,
103'h3b5b5d72822870174200000000,
103'h3f07150b5ebd5f12f700000000,
103'h1b0c1de3d918bc8578fffffff8,
103'h1e0e39b7d71fd190d600000000,
103'h1554b1f1732bef74ae00000000,
103'h0cc39a42503a292c847dddb76a,
103'h22efe1a6248edb1df600000000,
103'h1134e58f705275604671381795,
103'h1499bb09924257066a00000000,
103'h0d2a7ff862773c95dabfbffefd,
103'h12f56e13b610f79f6c00000000,
103'h3e4f374d023b7797cf00000000,
103'h18fb75e69730e5ab8600000000,
103'h06ea0b8694801cf88800000000,
103'h144fddbc6c7b92df1e00000000,
103'h1ac6a791b2659e65b200000031,
103'h2578e8fec8b57c222000000000,
103'h025c1017627c23b3d210176200,
103'h36bf542886f50cb29a00000000,
103'h169e2b18cb511cc9fe00000000,
103'h28e2a06ec01070f28400000000,
103'h04dc91e6d6ae9c0b4e00000000,
103'h0252a712be913c7a0ea9c4af80,
103'h06bdc8f1426dce60e400000000,
103'h167a0799c4c07573a400000000,
103'h2546b734cc7e3e64e600000000,
103'h0ac202db22f845feac00000184,
103'h2ece8afb873efd337800000000,
103'h1448e17cd101000e9a00000000,
103'h0083ad71becf8b0a20a99c3def,
103'h393cb7cb95186c86f200000000,
103'h12ee0824149c19f8b000000000,
103'h34de55b00ed8d1c44400000000,
103'h26cfa34aa0c6d9e85a00000000,
103'h16907bef54a52f986800000000,
103'h1c69c11afa74d2e30800000000,
103'h36df203f53054ed25e00000000,
103'h1f2d5127ee6f0fed5800000000,
103'h27425bf8e44e302caa00000000,
103'h04fc9662427b81549800000000,
103'h1e2ba3aea8bddd4d7c00000000,
103'h095fffcd6eba73afbef2c63168,
103'h23036bd98ce6175e6800000000,
103'h1ef508125546172bd600000000,
103'h1e62259fb74983056200000000,
103'h068d207a963e8b17b600000000,
103'h1d728f0534a0b0b76e00000000,
103'h3f3e14ee3b2dd1320500000000,
103'h354fb20316a060373800000000,
103'h22aad21d54de75257200000000,
103'h26447d4f492e27288800000000,
103'h1f7ed938acd8f945dc00000000,
103'h10e70654121d76952464c7df77,
103'h18ef93a6b29c4fcdd000000000,
103'h34d6961ec2835621e400000000,
103'h1aebbfbf5d72e9c896000ebbfb,
103'h2ad9e2a5d0497fe75800000000,
103'h0ee57c216a353fa6b4129e1010,
103'h248d656ad70f224c8600000000,
103'h3eb8a4d624f49e6df000000000,
103'h3356ce0a0a8203d8c700000000,
103'h393e7725493aa8aeec00000000,
103'h2a5b5fe73a9176b8f600000000,
103'h30876af5b4cfedde3e00000000,
103'h1ca814721e2b4dc57800000000,
103'h124ac1c74eb2b8bb2c00000000,
103'h112817cb6c5acd2d4a66a54f11,
103'h0a96e4887ea58ef49a00025b92,
103'h36d59f23d0cda6c00600000000,
103'h033fa7849a648b48847f4f0934,
103'h1c5c68a0903a2a6c5400000000,
103'h22d3f6e9d279d1f0ee00000000,
103'h26f11427aed63a918000000000,
103'h3cdbd82590aa317b5200000000,
103'h2b2b276bf89b45a30200000000,
103'h2ab4a11eb4771dc89200000000,
103'h3eb7ecc25ea245348b00000000,
103'h009172f78a56e6533e742ca564,
103'h13152aa8090ed3159e00000000,
103'h1f3427fb88a0460d2800000000,
103'h1cca43179ab570b53000000000,
103'h3a02a36838e998b0b800000000,
103'h2291ea0c16b3dbc85200000000,
103'h123003c590b67f308c00000000,
103'h0b6e638c3548693ca200005b98,
103'h1e62340806786d023200000000,
103'h2b3f9d3492e6d08e6600000000,
103'h0cd0e229714904966eecf35fbf,
103'h3f18a64eda88a1cb0100000000,
103'h26a8d3b0e75983f47000000000,
103'h14b16e1525722a434a00000000,
103'h14a0d907cb1afdf43000000000,
103'h04d94890decc6c095400000000,
103'h0e9a59e4f36d45112004208010,
103'h3eb4ef2d76468da1ff00000000,
103'h1241aeb944e0e786f200000000,
103'h32e96c394295d6b46900000000,
103'h335d95c296d7856daf00000000,
103'h243f045d08c0f1a6f000000000,
103'h0c6700997a1e8769863fc3fcff,
103'h3a6fe45cdf5d8bc69100000000,
103'h2d0e9ed4acc48c600a00000000,
103'h3284deba273470bceb00000000,
103'h02bc104693430f9196411a4800,
103'h0f11c93c86c7ee4bbc00e40442,
103'h38c50df90883fe925000000000,
103'h0e3cdf159695c7ced60a63824b,
103'h0ae920ef0e5ad5c7de0000e920,
103'h1ad8725a1c97b4dd760000000d,
103'h308fb210e880d5cc8400000000,
103'h10caf05a03594826a2b8d419b0,
103'h069bf671f4e8fa378a00000001,
103'h0ac7d251c4b3ea918c018fa4a3,
103'h2c8b630f0a4fe1038000000000,
103'h36cfc998d417b3554400000000,
103'h056d784942a316644e00000001,
103'h04f421313972dffd2400000000,
103'h0a2eb4aabce0584666000002eb,
103'h18b92927c2d479779e00000000,
103'h3d5b50fa0d032e225c00000000,
103'h22a08f30a4bc574a1e00000000,
103'h0358ad646317a8442a46200000,
103'h1ef123de84b83774ce00000000,
103'h3c5e13d04610e4d93000000000,
103'h26ce31e4650208b7b600000000,
103'h34faa742a0601c87fc00000000,
103'h263ec4e5072e4e6c6200000000,
103'h1d3b19fc3c28f5af0200000000,
103'h194853eca367ba940a00000000,
103'h3b579694bea2d4904600000000,
103'h3ec6f5c4d6eb287ce800000000,
103'h0964a3615342bf11a6130e387a,
103'h0f2b46acd009b4d67c04824228,
103'h3759a48c586e5837ce00000000,
103'h1d2ad6fc26999ee49e00000000,
103'h18e731e8dcf34370f600000000,
103'h28e64be7381e1a6d1c00000000,
103'h06ef1abc10054c55f800000000,
103'h3e6641c8b8eb983d3000000000,
103'h1b7707ba00dab2f942ddc1ee80,
103'h157b111c3e40f4c1fa00000000,
103'h049d34eb98b7fc7bfa00000001,
103'h06c4a510ec330d983800000000,
103'h02d7ad7372d04283d2ad737200,
103'h3cc568cf3894e794be00000000,
103'h36f418ecfa6c95083000000000,
103'h08dac586b931fdd76af59c28e9,
103'h06f47fb8ae2616c46400000000,
103'h38de7c6e7600dc4b1c00000000,
103'h225d60b8fcf55c03ca00000000,
103'h0648da0bb4d3d8724000000001,
103'h24665135d731392b3e00000000,
103'h2ea9df245e7a1336f200000000,
103'h30ee495e02e0646cca00000000,
103'h2e280f9b708a43912800000000,
103'h2035ae4b21788cef2a00000000,
103'h2a7486260ea09c8a9a00000000,
103'h132d7137f0d64ad5bc00000000,
103'h3cc6c0b69a4ad0fbca00000000,
103'h18ea53c66e784233ba00000000,
103'h148673c56b3f02ea5600000000,
103'h1ec3304f032956b0c400000000,
103'h1ad637ae56afca762e000000d6,
103'h313410097772fac53200000000,
103'h350a2a98504932738800000000,
103'h231f4811807d427cfe00000000,
103'h155dbc3b74876d154e00000000,
103'h1e4bfadb96a6b526ce00000000,
103'h1cad3440ec0471624200000000,
103'h2d57a019cb506c3dda00000000,
103'h3a7f4e6fa6fda07ec600000000,
103'h3e2e69dad35540989000000000,
103'h18843a6cced48f083600000000,
103'h1ede7c610d02f8e30a00000000,
103'h2e892a932487334fd800000000,
103'h253179440365afb0e400000000,
103'h2f2f088d70eeda440800000000,
103'h060126df152053880a00000001,
103'h2ad63e13c54f5c157a00000000,
103'h323288984a5082f48f00000000,
103'h3cf482cdb626c1085200000000,
103'h36a55747295949a09e00000000,
103'h07767f48a74dcc6e5400000000,
103'h1897035f9cf323b57c00000000,
103'h36080a6b2269a2fe2200000000,
103'h0a9fd27efd00a65dc04fe93f7e,
103'h0890e4337208b0c8e24c2a7dc8,
103'h2acfc2563ea88347de00000000,
103'h2b01c42e8739677b5200000000,
103'h0e9d6904f10929d19004948048,
103'h2d39b4391d0aee001600000000,
103'h3edeb0362aa857050700000000,
103'h0e2c2f7b16e20b3e2210059d01,
103'h24b3163b56c0bb744c00000000,
103'h2c4326cd24eceaef6400000000,
103'h0ede255f0aa0012aba40008505,
103'h1d217af5f6e327f7de00000000,
103'h0046dbcb04c14d56e8841490f6,
103'h3a2cf81460e2c84cde00000000,
103'h18ffff4d2129a417e400000000,
103'h027307b09a569c2c44e60f6134,
103'h20c9380bf5569b796600000000,
103'h04e0b5be36c9a32a0000000000,
103'h0adafbbd5692db35f40000001b,
103'h30fee5d45c7390f42a00000000,
103'h31796c17a74e8cb18200000000,
103'h274a8dd4574d7285de00000000,
103'h10e552bb06c6de9d840f3a0ec1,
103'h1212f2d7ad116c71da00000000,
103'h30b423e87ef6bf2ce000000000,
103'h34a3e1aad109b2048e00000000,
103'h0ee111f302bdd5ed0c5088f080,
103'h30e520d8b661b797dc00000000,
103'h3efa9c304642c98adf00000000,
103'h0b06d6b4b727ea639600106d6b,
103'h271cc33db5228693dc00000000,
103'h06f085b3bf295d489200000001,
103'h1c25ffc1a54620864600000000,
103'h389e435a6b36a63a0400000000,
103'h0a3e7156c65ca5fba8000001f3,
103'h100125e6fefae95614831e4875,
103'h14ed37bfc8395aacda00000000,
103'h3c1f6a1ed93a8093db00000000,
103'h108842b7ec27b853a230453225,
103'h2d4dc14cab4722727c00000000,
103'h060e29377acf652a6800000001,
103'h2807ebcf261d26771200000000,
103'h243c2efaad2b4fae8e00000000,
103'h0e982a79d6333b7db408153cca,
103'h203b486b7b6f6a786200000000,
103'h2eadcb87890794f23800000000,
103'h253d751aaa42dd5db200000000,
103'h06f86e5c58f0a8e53c00000000,
103'h3ee6a31bbd2e1dffe600000000,
103'h3044425382268c5c3e00000000,
103'h2ca9767d810d2f77fc00000000,
103'h13518805325171cb7e00000000,
103'h12ea42721efae8490000000000,
103'h0eb11adef34c704e3200082719,
103'h0c9e7fa80436b2c0505f7ff42a,
103'h0c9913e912e7cd9f427fefffa9,
103'h3ee519f59e864d474700000000,
103'h112c084b2c1f61305886538d6a,
103'h12bf66eeeb047b25f800000000,
103'h1a897852fb308371240000112f,
103'h333b57564eefea600f00000000,
103'h2b7383a0e97962b30a00000000,
103'h0ecb111bdab4ba0958400804ac,
103'h1f2719bcc7283daa4000000000,
103'h28b3a5ced4f34ec61a00000000,
103'h00301c40f21a6882e0254261e9,
103'h0025f5661ace0e51b67a01dbe8,
103'h1ad088949afe2a92a800000684,
103'h3ca3596d5b241ff8c500000000,
103'h3369790c36f4a88d5f00000000,
103'h1b4a012df29801fabafffffffd,
103'h1ef897a165017b06f000000000,
103'h3ea558a77f4b7c34e200000000,
103'h397639a65f4413d64600000000,
103'h293bc3329ce96c7dc400000000,
103'h0a994eb9945fa6242200002653,
103'h10f855477c9b6956be2e75f85f,
103'h14a2d80a4634b8105200000000,
103'h38916ea3562d0d57ce00000000,
103'h366971ba2acfe5621400000000,
103'h0aa11af5226154056a00000284,
103'h19742d86dacac5bf9600000000,
103'h2f7bf828e46be0b4b800000000,
103'h18b0d022bce00e3b9200000000,
103'h2eb58d7eaa5c06647600000000,
103'h291b9ee0050cd6873400000000,
103'h3a4c7600f2c26405de00000000,
103'h32e92dd69ade02e5e300000000,
103'h2765f3e7d72a78e6d600000000,
103'h053ec05d8813a6bd7000000001,
103'h2924635a6e799aa54600000000,
103'h3ecc6a5d32b85b02cf00000000,
103'h2e527445dadcbe5d3c00000000,
103'h3602f71558a928ba7000000000,
103'h04c720a248fb9d004a00000001,
103'h0304e4d47efe9415a4a8fc0000,
103'h32fb040982c5b4b7ed00000000,
103'h3ccde19bc4ca998c6a00000000,
103'h2049e7e876c59d95ec00000000,
103'h0cc18b3574937f31b269ff9afb,
103'h3637c29814dd671a2800000000,
103'h2573aeb2a29ef24f9c00000000,
103'h167a345998d6b4e7b200000000,
103'h3e4657967d4a639a5400000000,
103'h1ca5fa0512c497f3ec00000000,
103'h0ee3038dd30aef8a6a0101c421,
103'h22beff662eb0e98f7c00000000,
103'h0f71b0263c93ed1d4e08d00206,
103'h396ec4809e52ec837d00000000,
103'h363070ceecc49ca9b800000000,
103'h04fd0ca7a633612a5600000000,
103'h037a920fdd63d1f944f5241fb8,
103'h3a8c04956160dea0eb00000000,
103'h12f0639e62db70b0c600000000,
103'h17195f511e6775462600000000,
103'h0175bc2e3157d8e48a66ca895d,
103'h0735eb0487713835a800000001,
103'h2d56f87bc6e6f463d800000000,
103'h375376a3cd1cdf685e00000000,
103'h1eb76a11f973d7e42400000000,
103'h37733664b0c74e87f000000000,
103'h14a03aed0e7eb899e800000000,
103'h38b433d946f1eefe9900000000,
103'h28e50c2dda9229eba800000000,
103'h1289bc6695465dc4ee00000000,
103'h2af5bb273c2b69f2c800000000,
103'h12e07281ceb526595c00000000,
103'h00bd18dafaaae1809ab3fd2dca,
103'h0a2be91fcc8b5402680000015f,
103'h26e117298e486cdd6200000000,
103'h00c1af26197455fd301b0291a4,
103'h2a576d7bff556d26be00000000,
103'h0c980d5281171c4cd6cf8eaf6b,
103'h3d64012b6a6e89c8d400000000,
103'h3a7861e1b606971b5500000000,
103'h11011895346a9846be4b40273b,
103'h26df3c6f6ee2fa287600000000,
103'h3ad47c9680e412bdaa00000000,
103'h3b38468666c34f2d1800000000,
103'h30a2a791a097cbc39800000000,
103'h1a77a0e39ad01249fe00000000,
103'h322f945e0b72b9dba100000000,
103'h0ccb9a9624ea5abf3a75ed5f9f,
103'h0b2aeffb5919ef1d4612aeffb5,
103'h2b22112424e589b36a00000000,
103'h26e94496ee1079aec200000000,
103'h2d2331e55a328ad2e600000000,
103'h174779f3011bcf69d600000000,
103'h1a85b11ded3f014f3000000042,
103'h00a971fc42867b423097f69f39,
103'h16ddac895d0c2c601c00000000,
103'h074471e95eb59e5c5e00000000,
103'h36c706b334934ae5bc00000000,
103'h12889ccc3cd7bccf1a00000000,
103'h32d0ae27729ec3824f00000000,
103'h2f24ebe2c627604e8a00000000,
103'h092ec7fa78f80e75feeb64c7c3,
103'h16cbeef7e71cfa58c400000000,
103'h2340d2c46f4bc2533c00000000,
103'h20547a134517b14b2200000000,
103'h248f81b0a758840f9000000000,
103'h20c297c406acfe22d400000000,
103'h0212a8302b3c7fd37c40000000,
103'h12ae7aef8aff17978200000000,
103'h2661fefa0d11bfc7ae00000000,
103'h226e07141ec03ab73800000000,
103'h27270d51072239b14600000000,
103'h141c9361689040c56400000000,
103'h0c1131094eb74e166a5bbf8fb7,
103'h12178e78e2d3e177d400000000,
103'h38de269fb0e512812300000000,
103'h22c6f877c2fca0fa0600000000,
103'h36400b153adac799b600000000,
103'h1b706bc91ea1c01178fffffffb,
103'h2074adf4d4e1cb26b400000000,
103'h165e02a1af5236efd200000000,
103'h0e43f8488ec6e4e4a621702043,
103'h0204b5892524e78656d6249000,
103'h156732db3468dfcee400000000,
103'h3cab7b53f76d95580b00000000,
103'h1341fabc8cd4c8333e00000000,
103'h369f5f09c88043873400000000,
103'h0121aadd5ac23e43c0f1f4908d,
103'h3e0cd67fd0619d4d8800000000,
103'h3565977a5283482ae200000000,
103'h349320a810901eaab400000000,
103'h3e40ed5d04f5b6250600000000,
103'h20b0f855ba88d6cd1600000000,
103'h1482a09bf8c9c42a1c00000000,
103'h1ad7910d197abc7fd6000d7910,
103'h32bca028eefd5d1bcf00000000,
103'h0e976569c8d4ee28e64a321460,
103'h24fb0177ba918e51d400000000,
103'h322861afc928f3bb9f00000000,
103'h18d07e67ac23f5335800000000,
103'h2e75f83b5f4c56e32200000000,
103'h0cf06037f81cd54ace7e7abfff,
103'h24fc56866692cd862e00000000,
103'h0731409072832dbe2600000000,
103'h168a1fcdd77f84448c00000000,
103'h052f55ee5eb0c4d4fe00000001,
103'h2af16159b43ae4a2d400000000,
103'h37463a4b386a3a913200000000,
103'h351e40fae25b9beae600000000,
103'h0975cbef18a1d6361eea0eec83,
103'h3d7e1bb84cc017310000000000,
103'h22c150245435e3201800000000,
103'h026ebf2190b3fed86443200000,
103'h0377ca09b5754efcba40000000,
103'h1d22ab27f6e40e1e4a00000000,
103'h008da377385bd827fe74bdcf9b,
103'h3a2e7ee6947e834ff400000000,
103'h0683592e570c26c72e00000001,
103'h044d8272d03aa5adc200000000,
103'h3afbb9d596bdfedc1900000000,
103'h2905c9605d0b814eea00000000,
103'h2a8e5c3b16073b248000000000,
103'h052315dcfe0d0484dc00000001,
103'h2ef2752ca89b60bff200000000,
103'h2e7fd3586cbe769cf000000000,
103'h0c18b2d31ab0ebc99a5c7dedcd,
103'h3eb8cd724a30bf220700000000,
103'h3165ec96574971f52200000000,
103'h0aae6c7a55023f676c0000015c,
103'h10b562fb45682bfdc2a69b7ec1,
103'h326d4545ce1698781700000000,
103'h1f55e6b260cbfb735c00000000,
103'h2087fa14123940b92a00000000,
103'h38bc4cdd328f276b8a00000000,
103'h1458cba41317217f9e00000000,
103'h3e0be2e30ad36e5cd000000000,
103'h0a8af5955e2c3a00e2000022bd,
103'h29434900df381ce3ee00000000,
103'h388ac3d7e8c312794d00000000,
103'h1ae9602e90065b7a2a000003a5,
103'h091b6ae208911f5212c53ad80d,
103'h1679af96627a7f80a200000000,
103'h0110112eac95ea62aad2fdc8ab,
103'h15698540430f99f90e00000000,
103'h36c954cc031fab27ba00000000,
103'h22ba43a9d6893067fc00000000,
103'h3125b2084e528533fe00000000,
103'h2b270ac9710cc8ddd600000000,
103'h2737fd83a1327ae62400000000,
103'h25689b658b5985af9400000000,
103'h3b2269af709183333400000000,
103'h1e2ebd2d54fa1e98be00000000,
103'h3347d989111c88482f00000000,
103'h269370caee4b45758200000000,
103'h25388dbc62931efe9200000000,
103'h126f2de109268fc98200000000,
103'h169fec9e6f5f1d85e400000000,
103'h28ed33a400ce4b66ec00000000,
103'h2a85c01f166e38055a00000000,
103'h0eb16b98c15b6ba95c08b5c420,
103'h3c03a6dbeae12bc87300000000,
103'h16b4ffa4fa9297613200000000,
103'h3334a3d4f6963e3d1f00000000,
103'h2622800a4d4b3de21800000000,
103'h196bc7e9017fe1b70e00000000,
103'h36963b9026a261c15a00000000,
103'h0e5346987e0e29aa5a0100442d,
103'h1ca68fddf6a4653a8000000000,
103'h3845170584f7abd30100000000,
103'h13637fe4229e3bb0f600000000,
103'h15244a841ae352b67a00000000,
103'h14f33ece6c46d29a9c00000000,
103'h0a669853406b1d1eb600000006,
103'h04d19dab155e5bed2400000000,
103'h22dadeb3dec4f4406400000000,
103'h18c77273249691eb7a00000000,
103'h3cfad8cd0671709f5800000000,
103'h22995c459e38e3127c00000000,
103'h1c963bab5c33bbdf8200000000,
103'h35580f517ecd18252200000000,
103'h32b074e31b6353d07f00000000,
103'h347a4b140ebb6321fc00000000,
103'h167d0457816bd8051600000000,
103'h14b3797a76e623192400000000,
103'h10b706c28d632770a6a9efa8f3,
103'h271de7db2316a0eb1c00000000,
103'h0c402c15b2cda7ada866d7dedd,
103'h32ce48555aeb8f88cb00000000,
103'h0f4287ae272bbb9e7e8141c713,
103'h3719ee7798fa03f3d800000000,
103'h0307f62c273c8ba1fe80000000,
103'h00c3a58e5d567a19960d0fd3f9,
103'h186ae4795f5e7045bc00000000,
103'h163ddf02de2215d41800000000,
103'h2c0add80368cfa4d7800000000,
103'h2814679f8ccad9505600000000,
103'h00746bd878d5b6d08ea5115483,
103'h3832e05720ea1e701b00000000,
103'h11136aa9e35e8a4894da7030a7,
103'h1e80ef4a1a916a9fb400000000,
103'h38b94d3aaaa4d5499600000000,
103'h0cc761fbc925c493b2f3f2fdfd,
103'h02bf952d02df11ce5ca5a04000,
103'h181652a6cea673ca2600000000,
103'h0afe7ac0516608f728000007f3,
103'h288b78236a7c5b9df600000000,
103'h0e3e3a1a357ad65e481d090d00,
103'h36d00ddf5d064e81b200000000,
103'h2c08556eaa44889be600000000,
103'h34a6a5f52114967b4400000000,
103'h26c152198e1cebe9ee00000000,
103'h0e56d49c42c391df1021484e00,
103'h12f2a5a0aa84e3f89e00000000,
103'h00d2ff40f8dbb894e0d75beaec,
103'h10c7ef5c8ace5e358afcc89380,
103'h2ed9cb620aa15d768200000000,
103'h10af39469c694cd30c22f639c8,
103'h1a098b23cb4318351800004c59,
103'h1e3f9595daf2517bb400000000,
103'h2b43fe3d76fbdc9f7e00000000,
103'h02e9c45b953b72355a45b94000,
103'h36f8d74cbf7f7072d000000000,
103'h374b0273036934ce6400000000,
103'h108f7f14f8620c1b2216b97ceb,
103'h20cfd8566ead0e8e2400000000,
103'h044ba3cd3f3c8da31e00000000,
103'h2646dfb6de0c65f98c00000000,
103'h0cab506ee35809c6ccfdacf777,
103'h2b71cd420a9ee97daa00000000,
103'h36e558a3574a39ec8e00000000,
103'h029571a7c0bc072e988d3e0000,
103'h2e51f0a5b6a15fd1ee00000000,
103'h3d66796a7b36d179ae00000000,
103'h1519ebace888c21f6400000000,
103'h031797dbe4ef3b89def6f90000,
103'h30d14b3978092736c600000000,
103'h152c5e68fa20bf12aa00000000,
103'h34be43122af20a4c2200000000,
103'h3ad8e9dabe1e68b51d00000000,
103'h26e2cc2d32dcabc74600000000,
103'h08f5d5b66eb595a20620200a34,
103'h27299e52549861cf3800000000,
103'h2c4f713a5c8e3785a600000000,
103'h3293acd782b7d5d7fb00000000,
103'h2cb4943bf10747125800000000,
103'h128b1142629af3e9da00000000,
103'h0ef9f0180e4f8825ca24c00005,
103'h26f7067362da99682e00000000,
103'h00abf2a6b0d489803cc03e1376,
103'h0d6825ec56cb8ff39ef5d7ffef,
103'h3abf4d1bd677829a4f00000000,
103'h3665fc7122dfa886a400000000,
103'h16e7452e9c9ef5a27c00000000,
103'h253d176c5404f2139e00000000,
103'h0b5e799daaec37423c00000002,
103'h06f75e694f294eae9000000001,
103'h246febbb9887c84c3a00000000,
103'h20876eb05e7f26b58800000000,
103'h30a3e3b8c4ef12712200000000,
103'h2aac9003647681218000000000,
103'h34de8afc961a64da4400000000,
103'h16984e4200c6f4ddaa00000000,
103'h16d1383cf4a57fda4000000000,
103'h1cf934a90a3dce1c4000000000,
103'h0697b236a30f06593600000001,
103'h0750949e7e083b024000000000,
103'h06d06be4049fed38e200000000,
103'h3cf5c303caf081d76000000000,
103'h3e58e83fd0c0edbb6400000000,
103'h20cb13d50eb6b0bf2e00000000,
103'h03457a6c8d0f98ff00a2bd3646,
103'h265fce3cecdaacd40e00000000,
103'h166aa3e4af2027409a00000000,
103'h17366747d67ff57d8600000000,
103'h24b8db6a2cea99623600000000,
103'h3f4ae88b832100aa0d00000000,
103'h04b7a280e6d9dc143800000001,
103'h3b4483b6e524c49fbb00000000,
103'h06515a6a68dc6720a000000001,
103'h3f48ca802520ead78500000000,
103'h38613b3fea724541ed00000000,
103'h19538813eabb0fc21000000000,
103'h1c6a9987a31c4b01fc00000000,
103'h0b5e121bfd6fd315e6000015e1,
103'h1a727587d8da6c9d880393ac3e,
103'h16f91e35a2387eb98400000000,
103'h3d3ad6a57eaaf4415e00000000,
103'h0698da1754a412770000000001,
103'h0b66b09f12dee91c7e00000001,
103'h290ef3c45977c333d400000000,
103'h2aefb5a322de73d2e600000000,
103'h297b6bc34ced67973e00000000,
103'h3cab345a76dd1d3a6100000000,
103'h22b9e60e1e5888fdac00000000,
103'h21405af59c03bd582200000000,
103'h02a543affebda36642a543affe,
103'h2ef79401a0fdfe5bde00000000,
103'h1327018da2a3420bdc00000000,
103'h14aef817509ad60d7c00000000,
103'h323aabf922c1d79b1f00000000,
103'h0e8403413770cfb27000018018,
103'h0ccb58e528ab7bab9275bdf7dd,
103'h2ab5f094f92f7eecca00000000,
103'h1b3b5e5244fad7d1f2ffffffce,
103'h2e82a3aaaeb0c866ea00000000,
103'h393ab8b58aec26b92f00000000,
103'h2a9e496bf96eca63de00000000,
103'h1731590f30a983196800000000,
103'h04bf40845b47cc856000000000,
103'h22fdf060717925949000000000,
103'h0b28c6f5b6386618ea000004a3,
103'h2ac267eed93656795c00000000,
103'h3b058c01655f1d6f1200000000,
103'h26907c994e21855dea00000000,
103'h029492c5ca27115f4e24b17280,
103'h14d10f0b30b78df89e00000000,
103'h3f43e1c9f34c20be6800000000,
103'h0f15d1f7c71d2fc9988a80e0c0,
103'h2c094783856111938a00000000,
103'h1423ce6e9376e38b5000000000,
103'h2cf5e3523e802b0ed400000000,
103'h361418f452a3f97d6800000000,
103'h064f7e5ffe99dccfa600000001,
103'h1aebf55f34adf5c3fa00000003,
103'h02ff4fe9bafd7423f8d0000000,
103'h2a92d58316e969832e00000000,
103'h24ca5499d8e8b96ce800000000,
103'h1c9bb080427b8eeffe00000000,
103'h0a1b022aa745e389d80000d811,
103'h3497c7f904e1940a1a00000000,
103'h32fdf74a8efc9634c300000000,
103'h0a4ce00902945e2dc604ce0090,
103'h271757b7769255785400000000,
103'h2827b2efc0df35815800000000,
103'h2e19a23226f68d38ce00000000,
103'h020827a94e1e40288e09ea5380,
103'h1a8b0b4e3d37e25ab600000008,
103'h28a0446b80400a040400000000,
103'h3894b30a1acb15524300000000,
103'h2f7faee1856b59bdc200000000,
103'h3288eae17c000cc7dd00000000,
103'h34ca093c2a7fbba96000000000,
103'h364b319adc08a68adc00000000,
103'h14976f4bd2d2afc70600000000,
103'h344f06ba891de161e400000000,
103'h1206aaf11cb550adb600000000,
103'h193e0ad1120457683e00000000,
103'h3d7e113be50b02595c00000000,
103'h3290c76dbd490d2a6f00000000,
103'h32c15f017ac71e665300000000,
103'h0ea74742ec57e5d40e03a2a006,
103'h3c9186ec9e1944d58800000000,
103'h0e86c8efacc08c187640440412,
103'h1cc5181d285213051400000000,
103'h26ca85b0f6d8dbf4c200000000,
103'h1d27d918d49df411ea00000000,
103'h309e71563b6879c2e200000000,
103'h32d595ac169052dbb700000000,
103'h1e5ecd07072ec431f000000000,
103'h00c0e056bb0459de06e29d1a60,
103'h36c0e7b8586326e50c00000000,
103'h272968dcd824073bc600000000,
103'h2d223cdd0ee4eef41e00000000,
103'h3949d50f340e57d0f700000000,
103'h0175c71f603094ae04d32de6b2,
103'h1e04e014987a69bd3800000000,
103'h16b8004598f030dc9800000000,
103'h1b500f6ab8f510f132ffffffd4,
103'h14f67660cead1136ca00000000,
103'h2ccd7204e8fd20a18200000000,
103'h1e1ed7663cf397025000000000,
103'h2b606da42ac109073a00000000,
103'h2c9714d348dfe06d7600000000,
103'h3e7acd3932404e11a100000000,
103'h395ba640a0d762e4eb00000000,
103'h2f30164a5e52301e1c00000000,
103'h10c58f5b56add65ebc0bdc7e4d,
103'h3a3ae8d9c4ddeca91a00000000,
103'h16f09069d4a37c047000000000,
103'h147d9adecede64de3600000000,
103'h2f5cd571e6cef5480a00000000,
103'h20e9e663bb4c9026da00000000,
103'h1654e3fea8a96598c000000000,
103'h20635d9e08934bfc7a00000000,
103'h3a503c1b9ee82ffb2200000000,
103'h3b0c0fe1414b8d992c00000000,
103'h341473cdba9bc9b4ca00000000,
103'h18c63d52f6a7d9960a00000000,
103'h040b52d4aabc4d63c600000001,
103'h0e38985182828ab6bc00440840,
103'h1ab16b67868ddd8b6600000b16,
103'h20c6083256c675dcea00000000,
103'h1c827e933077e1447000000000,
103'h02fb4257d03de976c6ed095f40,
103'h2cf690d32cc06809f600000000,
103'h1e7fbcd9eebbaa61c600000000,
103'h24cf5ebd9cb23b34f200000000,
103'h1c96e1e5bb31f80ee200000000,
103'h229c4e849f0156cc7e00000000,
103'h1662232d7a9838b23800000000,
103'h38e3a2381e348736d600000000,
103'h37175c77b496aa645200000000,
103'h2f7d0ec62d7a4c9c7000000000,
103'h04e417e12291a9142400000000,
103'h16e359ae510eb7da5000000000,
103'h061722b254f2cfbb7200000001,
103'h2ae1961aacd62969c200000000,
103'h3a26561f72ed4c1c1600000000,
103'h2cfcbf385ecee236c200000000,
103'h2ee1e02b98f538563600000000,
103'h06b9d0da46f1f78e9400000001,
103'h0867eaf2b4d3d7ba2c5a1ea44c,
103'h3e0351273a8da8947200000000,
103'h136d999284f593872800000000,
103'h00cd1a5402f8e4ae62e2ff8132,
103'h331e92a416667e40e700000000,
103'h1b43e2ae57339894eafffffd0f,
103'h3ef6db4d09522b390000000000,
103'h249f6772e4960de75600000000,
103'h0f40d847228ce9345e00640201,
103'h0e48c75c462c50a74204200221,
103'h24844f06566d28ee6400000000,
103'h041201e964b5f04aac00000001,
103'h0735c2b3cb3a3f510200000001,
103'h2ce66cb28e4c413a6600000000,
103'h18c36758948203ee3000000000,
103'h1a0d8aed006870a0be00000000,
103'h000d9ecc192bd7f9549cbb62b6,
103'h3247f1fc323962e65500000000,
103'h30ce8666b54701b26e00000000,
103'h04d71ebf668ef3aea000000000,
103'h1a4827b8d65d7a1554000904f7,
103'h08e508ab9c3498d4ba68c83f93,
103'h28bb4c84b77cc08d9200000000,
103'h3ed892103f61c9392e00000000,
103'h3884cb4a671d15bde400000000,
103'h0a8e7e99e4f5a7ce220000239f,
103'h38cccabe1e7a73188800000000,
103'h1c87d76fe908f1b26e00000000,
103'h3ea4ad5ae2d5bc708c00000000,
103'h08de9903be5d93e074418571e5,
103'h370e2c7abe02413b5600000000,
103'h02b8330a46e0da3f16cc291800,
103'h376b2b4c3cef06b9d400000000,
103'h0ef3dffebea739c41a518ce20d,
103'h24da2891b51265105600000000,
103'h38c2b2600306450f1400000000,
103'h128c166d66e06da0c800000000,
103'h284481349ea32000cc00000000,
103'h3ca425bff02f366e3200000000,
103'h04162f5b9973b7a2d200000000,
103'h108e7e065417dd62c23b5051c9,
103'h04e73a51db2e0cbe5c00000000,
103'h16e3169e2abc8ac4b000000000,
103'h180e2958aea3c5168a00000000,
103'h34acf3b60486dbb4b600000000,
103'h27639b761e95050d6400000000,
103'h30484ff49341f8c36a00000000,
103'h26e98f37b8a594398800000000,
103'h0d2e93916aede42e1af7fbdfbd,
103'h36fa739fd0d77365d400000000,
103'h3e5b58bb9d0606f73e00000000,
103'h18fe369ad2007a970e00000000,
103'h2c46a8b3915bd352ac00000000,
103'h2b7cfefa6a5a09ed7e00000000,
103'h3a8ac8a716a0b2a11000000000,
103'h269e994b031db19b7a00000000,
103'h24b2e485fca87a429000000000,
103'h35230313a247138d9200000000,
103'h2eed2b8ec6f9f8138e00000000,
103'h015806aafc1cfb2730ba80e916,
103'h12e09362ab0a26b5f800000000,
103'h22119a5ceb622d60f400000000,
103'h1289b4e4be42c0c39e00000000,
103'h0afbc78021545b208a03ef1e00,
103'h3e8ad542b2de10054800000000,
103'h1f2409bb3ed9d7856800000000,
103'h281f6b94bc64acc81a00000000,
103'h305d8e31da88b6835800000000,
103'h18f00bef82a822181600000000,
103'h326099b27205b049f100000000,
103'h0caafefacaf5bc39747fff7dff,
103'h235a110b3e5655ebe600000000,
103'h1291d99f0b0154e6b200000000,
103'h0771c44aed5b65f1f000000000,
103'h2e575f40beed3f90fa00000000,
103'h2132b670075f03dbe600000000,
103'h1164638b34b6631ca457003748,
103'h0a97658d14e9198caa0000025d,
103'h3125cd80e44d7d17de00000000,
103'h14a17505aee4e2a4f200000000,
103'h017c20665e0ab025d6c368461a,
103'h1e0d2ee3b2ac252b8400000000,
103'h128756edb2284591e200000000,
103'h294efc0f933574759600000000,
103'h2efb83d664bccb634800000000,
103'h10b2bbc30c0bc772da537a2819,
103'h261618db3a074b493e00000000,
103'h30a1bb854cba070c4c00000000,
103'h0a62d2a4f2d01fe786062d2a4f,
103'h0ae0b527e271db6cd200382d49,
103'h176a5f1daed4ae11c600000000,
103'h1cfb545cb8b56339a800000000,
103'h314650a80e1fc2575600000000,
103'h36616cdaea1b16b40e00000000,
103'h1eee647a9a61675c1c00000000,
103'h36500a2c10c2d4370800000000,
103'h0567131730b138b1a200000001,
103'h229dde59a70142ddb400000000,
103'h2aefc0502b6855f4e400000000,
103'h0ca309a2cd06344e8ad39ef767,
103'h0019272c76f5f49eb4878de595,
103'h25407d67c498fe418200000000,
103'h2e691680c4b2256df800000000,
103'h24fa058eaaf2a2d5bc00000000,
103'h269128eb195bb9568200000000,
103'h1e1e40e63d55bee52c00000000,
103'h1c445722e2e6e7d04400000000,
103'h1f1c92cd830528b68200000000,
103'h0ae7714dde497fd96400001cee,
103'h0f0e0924bc6612a6e603001252,
103'h108a5fe0c64d83f4c41e6df601,
103'h36ed9e6d145b8d198000000000,
103'h1d5605afe6e5ecfa4600000000,
103'h2307eccc1cd38b675c00000000,
103'h221fe68f392991174200000000,
103'h2a8564471b317de35e00000000,
103'h07466f187e5164729600000000,
103'h08ed66e428d6c8b9b21dd72ecd,
103'h2767ea172f1d37d23000000000,
103'h3d0bfe61770a9eb65800000000,
103'h2ee1908f1d7288cd8600000000,
103'h1e08872f597e872efc00000000,
103'h37064689496017be1800000000,
103'h3c213db566689eed7100000000,
103'h3946d397de6ee576b900000000,
103'h10def247da90232c2027678ddd,
103'h02f59826d4d6f6c3fe00000000,
103'h3a6c55c3e4b5e90bd800000000,
103'h1a4bb24e66ab8132ac00000097,
103'h1899f44fa317d6f69200000000,
103'h3278597cfc638944f900000000,
103'h1f2db56e56fd7d949a00000000,
103'h3098fa6b8975d7119800000000,
103'h2aafc09b66a38c7fee00000000,
103'h04de5dc1d93c86eb7600000000,
103'h1d70842d42ec4786dc00000000,
103'h0a00282d46caa548b400000000,
103'h0105a33ee43b2975f6a0665a6d,
103'h1eaeaad06f3b51a33e00000000,
103'h1294394d7140f4e22200000000,
103'h0b660f514eef9fb29000b307a8,
103'h08028a9de083d9000040a9cef0,
103'h2ada2f606ae9e8514e00000000,
103'h3aed25c632ec72ef3100000000,
103'h3c41110e1cc6a24f9b00000000,
103'h0a849c0898b3c815ce00849c08,
103'h3b4c000314f4d923ea00000000,
103'h16fd4c4ede79752c8200000000,
103'h249b0b89dac5752f9600000000,
103'h0eff6d1470c2c17e7661208a38,
103'h131796b4d55dcd085000000000,
103'h28249979235d3a1cc000000000,
103'h1eab1169f574d0d19400000000,
103'h2ef6fe8a5e996a4ab600000000,
103'h2e05ad293d447bb4ac00000000,
103'h037228d06d3b7a3f0a228d06c0,
103'h3a3bde945a4127684600000000,
103'h277a6529deb35038b200000000,
103'h3152560a18ef2ecd0e00000000,
103'h376ec29eff6993f6ec00000000,
103'h2ac6a972eebbea010400000000,
103'h385fb7af252aaca00200000000,
103'h24ac16240ef15612f000000000,
103'h28e7a36606510dc21400000000,
103'h2a8cc49eeafd23e62400000000,
103'h1aedcfd8d2e4c74c2a000003b7,
103'h2e7987b2bd718beb1600000000,
103'h12f6959f965f5bc3e800000000,
103'h3ec4b14e86d8e376a600000000,
103'h148ff0e398cf79163c00000000,
103'h3c3ff7c4d6942a64c300000000,
103'h22618a912b241b485c00000000,
103'h20e279216864130d3200000000,
103'h223c4b284ac59d9e5e00000000,
103'h3e6596456aa816bfc600000000,
103'h33230bc74ee461e81100000000,
103'h10049c918d49f82d7c5d523208,
103'h164a4068ff6d03f4ca00000000,
103'h265581dece71a0865600000000,
103'h2208da1464bbe0ef5600000000,
103'h2ca094320c1162ce2400000000,
103'h0482467d2f1a3ce28a00000000,
103'h1ad0fcbd1cbad11496000d0fcb,
103'h3e915383603d1791c500000000,
103'h090d8b38fa0e144ee081cfbb0d,
103'h1e9b25bcb89f67d24000000000,
103'h2542fd2302acf30b3a00000000,
103'h04a5a59de14818c7f400000000,
103'h064565aa848b15eaf600000001,
103'h00f33a060a30bb88d691fac770,
103'h35407633d17621335c00000000,
103'h2a3aa56cd1695b396600000000,
103'h037ced6dc6a9d16d3618000000,
103'h1e4a4b59b0e476da0600000000,
103'h044864ce72616447cc00000001,
103'h3abc9f7690abafa17f00000000,
103'h009a355814f4146ff0c724e402,
103'h0e219ca6ceb0b3e68210485341,
103'h0c8d7acf904ae93e9667fdffcb,
103'h3d5abd401f6c85e56700000000,
103'h3ed3af522afa00b4f600000000,
103'h1640b5d42754bdf51400000000,
103'h3d5e703ca7286d473e00000000,
103'h32c713e3bc69231b6500000000,
103'h069c3d7038c793580a00000001,
103'h056b67b1aa8ea73bc600000001,
103'h288f4fe8302ae4abfe00000000,
103'h34dba565f4964c5da800000000,
103'h3a911dff1c259c45d900000000,
103'h3a0e29f0500141abcd00000000,
103'h2319dd1d4c925faaea00000000,
103'h3d5074f646a0899b3a00000000,
103'h081d592ce8ba66b886539fca37,
103'h320fd9a9640adbaecd00000000,
103'h2f039bd1af2834dbb600000000,
103'h3489bda4e0380e851a00000000,
103'h02b069134e3baa56c883489a70,
103'h38917b3a44c567fbab00000000,
103'h137d69100675d10ef800000000,
103'h1c918bc17e074c493c00000000,
103'h06ddbcf81084b5594200000000,
103'h3e6598856c16411ac100000000,
103'h3cb2dc0e72f3fe12d300000000,
103'h3f75f0a6725996983f00000000,
103'h01405187af0c72a6b226621730,
103'h128f67c22c82634d2400000000,
103'h10f4bf176cc2b4d4d21905214d,
103'h024e147f7e521c96fe80000000,
103'h2701007fd146dbae6c00000000,
103'h38c05f26d294f02dea00000000,
103'h3902211afa95f0adbb00000000,
103'h240697e3f3564fd48e00000000,
103'h0e5d2b43eb5870ef882c1021c4,
103'h0afa9a524e5f08d37a00000003,
103'h192cf98e9ebc34176600000000,
103'h20f54978a8b6ce69b400000000,
103'h1b13e93740e3c7f852ffc4fa4d,
103'h008af9e560d91170fab205ab2d,
103'h36611366faecfaa83a00000000,
103'h08f360fffc77f48d9a424a3933,
103'h053c7d02b2d907f49600000001,
103'h3e6960fdbacc68f49200000000,
103'h1a6f5669bf08e5f7440deacd37,
103'h3162467dfe7246f4fe00000000,
103'h02cd2b1fd8e19d5ebe00000000,
103'h071117b64943e3dcbc00000001,
103'h05216d414b110efc9400000000,
103'h033aa8c3912226b2dc18720000,
103'h3ec62b3ad54393f42600000000,
103'h13334b10d97e3cb7b600000000,
103'h2ee44ec3964467f28a00000000,
103'h14a66172ea77b3036200000000,
103'h0a8a9ad5195c01c6fa00000002,
103'h16b2682b6f026339e400000000,
103'h38587239788cfe0efd00000000,
103'h3242e43a0e3f663a6b00000000,
103'h16a5093e0897d873e400000000,
103'h14633008fadabcadf200000000,
103'h3f23ba0dd27fc5ebfb00000000,
103'h23714221a6e2f5f4f600000000,
103'h16fe306fe506b002c800000000,
103'h1122f7320977f2246ed58286cd,
103'h07227aa21e7622945200000000,
103'h0ea1c3fe2e9919c65a4080e305,
103'h3d04034f36bb94687800000000,
103'h106cf2a3055d5866a887cd1e2e,
103'h2b4dd41b43615bb5de00000000,
103'h24a4d827d2ce4e58e200000000,
103'h0c94f5fabc1c2274244e7bff5e,
103'h2a40a83620c0fa9bf600000000,
103'h0c49b2d82d55f096b4aef96f5e,
103'h32b41930169698ccd500000000,
103'h28eccde0e4e04ba50200000000,
103'h1d41a505d69464d51800000000,
103'h325776c6be8132b5fd00000000,
103'h34c3391e5cc2d7bbd200000000,
103'h0cc59442cf1a4e8292efef616f,
103'h0aa83b0c42dd87a0ee000000a8,
103'h1c1f46aacea31be3bc00000000,
103'h2e1784ff594b56effe00000000,
103'h1cd29b0fb66a9d9acc00000000,
103'h18a7ffa2a482229a2600000000,
103'h175aebd68354bda9dc00000000,
103'h24b0f3ee1afcbd4c8000000000,
103'h0b5252f5b257a923025494bd6c,
103'h275e4f9817089d111e00000000,
103'h26ec6ed4a15af006d000000000,
103'h2acf4bbb06b93f9ee600000000,
103'h08aee5edeca5ae738605a5cf35,
103'h18e62943d774fa2e8c00000000,
103'h3e2609aade23e01c7900000000,
103'h04c0da18b70a09605000000000,
103'h1014ea257430130b2ef26b8d23,
103'h080ea8a5b8f0ed23e67f22c32f,
103'h187d61548805d7495a00000000,
103'h090ffa1fd3147fef140dc2f863,
103'h2eac9c4b6a91e1439c00000000,
103'h0879518232a1db636e6c4570ae,
103'h1c36f3dce14e77aeda00000000,
103'h3afa6d80eac7c9310d00000000,
103'h28d2671406febd0dee00000000,
103'h023c41eac0f92a8ed80f560000,
103'h1147f824eacb91a2de3e334106,
103'h3ea2260ded07d38da000000000,
103'h16c41d27fd4fcbb28a00000000,
103'h34e4d14ffaf1f1c07600000000,
103'h14feb006d0b60ee87400000000,
103'h1ee42060869ae0386e00000000,
103'h16d16447da99903f4000000000,
103'h0b0e73e1bb7db09fc610e73e1b,
103'h393d753c104f14e7a100000000,
103'h3922857eda5d88c95b00000000,
103'h3ea275fa129afe056b00000000,
103'h20bbf6b48cbd83844400000000,
103'h3a53280ecb5ff97e5900000000,
103'h26396e50ab1bf032e400000000,
103'h2b7d3d5be66f1841ae00000000,
103'h035c0a6c8ca886925aa6c8c000,
103'h26f85b017725c3ee4000000000,
103'h16f4a514ba81ce5acc00000000,
103'h300cdf5ae07a295c4200000000,
103'h309431e2b66ece70fc00000000,
103'h3cc40afce77badcbdf00000000,
103'h3e19a805560fdfae9500000000,
103'h3cf1136892d3eaab7c00000000,
103'h1b42a82812ed92b0d2ffd0aa0a,
103'h2f030b588edea6196600000000,
103'h2b3f1c54e9214e417800000000,
103'h3e8b0cffd724599a0600000000,
103'h24aae856436375eeee00000000,
103'h1cb8565d80ee82eec400000000,
103'h22a46a7e24996b450600000000,
103'h10b1cce04051c1a28630059edd,
103'h14e388dc62f62c20aa00000000,
103'h1d78bac772a7f900ea00000000,
103'h22fc6fa1468b81dd4c00000000,
103'h0e198fc022043ca4be00064011,
103'h388871818700ac460600000000,
103'h06ed7f63941a3c062800000000,
103'h04fa86468ca2ad87ae00000000,
103'h0a930f06d2902ceb4224c3c1b4,
103'h352fd46bd88ab331d000000000,
103'h22cd4616e21dc238a200000000,
103'h2684f3c8164d96a47a00000000,
103'h36df4f00fb1adcbb5e00000000,
103'h18c9d725209fd0837400000000,
103'h153f127b167f1f846e00000000,
103'h32d21009ae48f6a98f00000000,
103'h26b2a43cc2880924a400000000,
103'h16ae152b355a192e5400000000,
103'h2549569d1c0cbd6b1600000000,
103'h0b63b79372bad2964c02c76f26,
103'h1ec70f33570429336800000000,
103'h34b26ff7e167e0c6da00000000,
103'h00f7e9eabe2eeffa30936cf277,
103'h294a2148b4e15ff21200000000,
103'h02572b3cf4d949dcd0959e7a00,
103'h35685e649e236b258400000000,
103'h06e17253217a96627a00000001,
103'h1689763bd4e2f4c71800000000,
103'h1c12da169ac4671a3800000000,
103'h177587ce334ddd560e00000000,
103'h2efba0ab4e60b76ca800000000,
103'h26fc4feae4d63f3ada00000000,
103'h34dff3f192d1dfe62800000000,
103'h1e87ff1278ce2fd10c00000000,
103'h397de7896eae23c29f00000000,
103'h22d4876d0d3622d51800000000,
103'h2e01668b84b40a5e8600000000,
103'h0e002590268891cb920000c001,
103'h26cd1465d689f8571600000000,
103'h2d4826fe248a1de73e00000000,
103'h3ef95c6b8b57324d1400000000,
103'h155e9c37769f594b3800000000,
103'h134c6dcef498b5b6c200000000,
103'h26c437bd88f751ee3800000000,
103'h1ec61f935d43bfbd2c00000000,
103'h201f39b64207f77ab400000000,
103'h1917ad2462ce170e1000000000,
103'h04a8d64942ed50c45400000001,
103'h3b31515c5d04fde8b700000000,
103'h0afd8c2ca0add431f800000007,
103'h1ed1be779adf258e5400000000,
103'h157407d0a6dcb1baf600000000,
103'h0e03a1ee04ae70329001101100,
103'h229839f41a2278033600000000,
103'h18daa62c292619f13c00000000,
103'h2afc37f28abe53e55600000000,
103'h20fa7b73e498fa117e00000000,
103'h1ca72f27ce9532040800000000,
103'h32765adeee8fad77ed00000000,
103'h316ba0874c36dc9fba00000000,
103'h3a1f3a14fead377eaa00000000,
103'h276bcdb43118d805f600000000,
103'h234d93576a38121af400000000,
103'h0cbf067290a3dfcf245fefffda,
103'h0267562d72f173268ed58b5c80,
103'h36bcdd66feb079992000000000,
103'h1c2b3ca68017cfc69200000000,
103'h2ad1ae00f8d4ad2d9200000000,
103'h0b1bff2a94ffe9d4120046ffca,
103'h1e57c37abed197d50a00000000,
103'h314401640aed96ff9e00000000,
103'h03480f13e9455a7a5ec4fa0000,
103'h0f20c9f158895bde680024e824,
103'h2cf96ea2dad16af25000000000,
103'h0aa3ab2968f234e3a80000051d,
103'h333b7eaf96eba3868300000000,
103'h0218acb0208f4eafec04000000,
103'h2b7f368f14cacd5f8200000000,
103'h2eb72b6056e37a0fa200000000,
103'h1ae155154262b09eb60000000e,
103'h1cf72250b119dbff0e00000000,
103'h3e9c3e3c0afb31145000000000,
103'h370c2786e6f253650000000000,
103'h045f8ae1648e91a10a00000001,
103'h14159eda9a9ab927f000000000,
103'h14e58ed2defa44095400000000,
103'h1eb0afdf730fe2e3f000000000,
103'h0e6e245106f571b6ce32100803,
103'h22ba2a63a4a621964200000000,
103'h12a0e99e321445e74800000000,
103'h2281ece216ce704aee00000000,
103'h2472d309e86f59e92000000000,
103'h2c592ae88af146cb3600000000,
103'h1ae5a45d6f6419d520000072d2,
103'h3c8663b99cbd44bdab00000000,
103'h32f59360b6a2e91b1b00000000,
103'h12d41cf0f3294cd4b600000000,
103'h3ea3ed4c661ee0356d00000000,
103'h18d7d77cf8f2fd266000000000,
103'h0ec9066b3696ea72c640013103,
103'h3a5d1e748e6ec1efbe00000000,
103'h1a1a83529d37c85af600000001,
103'h20f6c8661894e6cf8400000000,
103'h20c60a9ff2af6a222200000000,
103'h172c374c94a632883a00000000,
103'h1b0125e8f46c3d282cfffffe02,
103'h3d0ddce04a987474c000000000,
103'h36af7aa724999a5db400000000,
103'h2500829022a7773dfe00000000,
103'h24f7bd015956f1e52400000000,
103'h1a5b349abd5774754605b349ab,
103'h195720a8e24f31769e00000000,
103'h3ceca714bcaa66115c00000000,
103'h0229a4be950186ba3e00000000,
103'h22bd944d92ee2dcefa00000000,
103'h3ea8f851d417d28d8f00000000,
103'h3ce38dccb6d566db2000000000,
103'h36c88958f57e5f2cf600000000,
103'h04af0b9f7061ecf9ac00000000,
103'h2683bbb4e72a7652a200000000,
103'h1d703e57ecd981f21200000000,
103'h093227d6135d3da6fa378d3874,
103'h2b7270812ecd7bfee600000000,
103'h3e14a625f6ffa3d4f800000000,
103'h38e1521d637214562600000000,
103'h1e878006e086ba7c1c00000000,
103'h168aeb9758680c997e00000000,
103'h3d5bd326b6ef8ca05e00000000,
103'h192c5e8b0c7a7837b600000000,
103'h196efe4588d64b5e6c00000000,
103'h3638587c2002a9e97800000000,
103'h2e69bf4c3871a82f0000000000,
103'h1a8ab2bcb0aa00ab22000022ac,
103'h15261e64de13bff75a00000000,
103'h1497d56b789e72b40a00000000,
103'h360c365b8cc49118e800000000,
103'h12f23f7aa35c66846200000000,
103'h1c824944d8689cdfee00000000,
103'h062613066a5adc5a9000000001,
103'h29684f7c08dd259f6a00000000,
103'h176f1d0a8e0338a5d400000000,
103'h28d2511d766b8821dc00000000,
103'h129e22104cdaa52c6a00000000,
103'h26c4cf5db4acf649e000000000,
103'h04c8a24a874b185a2e00000000,
103'h2ecfaddd2e0fe7b7e200000000,
103'h11424191b2d88a026a34dbc7a4,
103'h3e8f7a72a0a837df9800000000,
103'h2089a99d70ea79714a00000000,
103'h0acef1226e79f3e3ea0000033b,
103'h2324205f51039d815c00000000,
103'h2c51d99e9ad28ea3ca00000000,
103'h1927cabd7ef6af031a00000000,
103'h34e8354dab4888a1b600000000,
103'h3e2293c1c370535f3400000000,
103'h1a608fb7365888acde0000608f,
103'h11711a50777b1c6ea2fafef0ea,
103'h057853ecd0dbac25d800000001,
103'h22c8162ae04cc6764e00000000,
103'h04882bc824c51a631e00000001,
103'h1ea0ca12468d308dfe00000000,
103'h2d3484cb0c155c562200000000,
103'h0ca3eba9aab626686a5bf7f4f5,
103'h0a6018fe96eaab337600000006,
103'h2ee160b6a28e96dd2000000000,
103'h18efd8fcaeeeafdbb600000000,
103'h0f13ad98dcd010925a0800482c,
103'h2eeda89d74bfe98f0800000000,
103'h24b24ed582d39727e400000000,
103'h3f058beab0c13fc55900000000,
103'h064778db95738e9ada00000001,
103'h2b59765ed5791a858a00000000,
103'h022b5d711ac093611e5c468000,
103'h1cd0dbab461a09bff200000000,
103'h263799aac94567310e00000000,
103'h0711e645271642dc5400000001,
103'h38654d650c4ddc871c00000000,
103'h067947e6125fc2cc4200000000,
103'h1aa74c270cc51031500053a613,
103'h381ab799123e58176300000000,
103'h3aa465e76ee5a43e6e00000000,
103'h0b7bf0bce7005bd7825efc2f39,
103'h2eb33e5ea0a4c1bef000000000,
103'h1caf9c31ad20b27bd600000000,
103'h1eea521c1ad3f0da7600000000,
103'h0e0aac44f6838d0c2201460211,
103'h252b6245566ddf283c00000000,
103'h1cf0da04a5788b6d3400000000,
103'h3ed7043fcaa3edb28b00000000,
103'h3c911f556694c7b72f00000000,
103'h30cec777246bcbf6f800000000,
103'h3a7a4ec120fceb4c5e00000000,
103'h289e617850cbb2c38400000000,
103'h226661e20a460184a400000000,
103'h00c32a02f4e462fcf6d3c67ff5,
103'h048bbe1ad64ac4df0000000000,
103'h2a513d7f160deee1f400000000,
103'h20e26fa6dc99acfcca00000000,
103'h20b9a35346eaea7be200000000,
103'h177539fca6cd5a22be00000000,
103'h207b95850686fd760400000000,
103'h028fdfef5cfc3772aaf5c00000,
103'h013dd7567e77ccf7b0dad22717,
103'h04d6b9398107ace70e00000000,
103'h2f3cf53f4345843d8c00000000,
103'h202a2ebb061c3d770c00000000,
103'h2f139fa9765932b64e00000000,
103'h3b74dd8f968361715600000000,
103'h06ddc85cc497011acc00000000,
103'h168c37677f0bdeaa6200000000,
103'h2c56e3e944e9a7072600000000,
103'h387ac3215b75de6ea400000000,
103'h1a2203cac6ccc257e800000110,
103'h0060458eff47857944d3e58421,
103'h24aa65fd986989440a00000000,
103'h0cde2d7358c9ced30a6ff7f9ad,
103'h1087d357bc7434d0a209cf438d,
103'h1cfe3b940b526243fc00000000,
103'h26bc29499ada359bb800000000,
103'h08e3a04336d8712fc21de8b67a,
103'h04d4e60fdc949a795e00000000,
103'h3f3a60ad26783abc9500000000,
103'h00f23d8e6b4d20cc721faf2d6e,
103'h1e84500b688781799800000000,
103'h34eed3b82a79bf080200000000,
103'h26edf1de48fe0f136c00000000,
103'h3e654ac0fcece2cb9600000000,
103'h0029c47022dad4a9de824c8d00,
103'h2c75bf98e1401f6adc00000000,
103'h033b79c9a269e3dafe80000000,
103'h22ff430dcedfa373e000000000,
103'h3eafef1d931b1d3d8200000000,
103'h3d3b6fd7341a604b5000000000,
103'h1d070ffbb2ca4f68e200000000,
103'h1e3c93fb2e05bf401600000000,
103'h3151bb6e8c0ccf3bc800000000,
103'h1282001f6b496336f800000000,
103'h2acca51b9a9b1ea58400000000,
103'h32e19980ae1d1ec4ef00000000,
103'h2afc4d25d8e9c3e08a00000000,
103'h2e23d006cacb5d613800000000,
103'h1e94b61eb6c7aa871000000000,
103'h28a0badc24eb7a8dda00000000,
103'h20c9de5e828030ac9000000000,
103'h30dcc5c16b20eb88b600000000,
103'h0abb0a858aeac9e73800000005,
103'h1c60f9d0bac78fa8a400000000,
103'h12f263a9c6829a2e2e00000000,
103'h0b03fe2f62e393feea0000040f,
103'h2f36843db4d5f7a8b000000000,
103'h1e53d4333ed9f5d81200000000,
103'h0938b3d16f107a15c61464e254,
103'h38a02d9dcc644e490400000000,
103'h0aeb3b69149d021a720000003a,
103'h110c40dd0c3d2fb83e67889267,
103'h15073c2916286b215200000000,
103'h0912b18ae634abfe5e930d3a5c,
103'h06827535ba3be8277400000000,
103'h1a8f3afb024e99b25a00023ceb,
103'h38d930788ad10ee81600000000,
103'h2f4b9117646049e31800000000,
103'h08f29db49c397a5ba265f3f79f,
103'h1ed592794a850b730600000000,
103'h390720f05577a927a500000000,
103'h1a09be4f724d3ba0ee00000009,
103'h226ca591aa545c914200000000,
103'h0709072f875e1ae0b600000001,
103'h352a744068cac0726000000000,
103'h38c38a78eed3c7a1e700000000,
103'h2ea9dc5262fe3be24e00000000,
103'h0ee48abd1ac1c65b3c60410c8c,
103'h367d5408896ba2ada000000000,
103'h04e0ddc658502d6aba00000000,
103'h03182f260ecd817344305e4c1c,
103'h224dbc6812ae5f399c00000000,
103'h1c45100554c68e5faa00000000,
103'h20a8065036144ac7bc00000000,
103'h3d5b2a05d5595acd1200000000,
103'h26dbcf2eb401611d4800000000,
103'h250ad391325c8b231c00000000,
103'h3600665359385a51d200000000,
103'h3e0a43dd3d432de30400000000,
103'h1c6d7c34324394365c00000000,
103'h2ed215a8734dd8139a00000000,
103'h32933a3fcebb5447cd00000000,
103'h0e8cb928fc8d69f03e4614901e,
103'h28c965f52e20a4300c00000000,
103'h3649a6f7bcad5d590800000000,
103'h3517c00de676c34e3600000000,
103'h02a12d6bdcc06a45f4b8000000,
103'h0ab804ba10d82a53da0002e012,
103'h02ef8038537957bfb648000000,
103'h36d4590f9e315c79c600000000,
103'h112ff5352120dcb21a078c4183,
103'h074bfba096f535c1b800000000,
103'h0d402c5fe7252af6d8b2977fff,
103'h26adb4deed7126976e00000000,
103'h1e4c99d7b8b152f75400000000,
103'h370c5b82a15f07d64000000000,
103'h24c152ef3eaba1adf800000000,
103'h389b7552b6b7fd309900000000,
103'h38e6be4d9b79501fd800000000,
103'h32e35a3fd514c5728f00000000,
103'h0a3efe084cfb83c028000001f7,
103'h2246437ebededdfffc00000000,
103'h31058625cb1ddc084a00000000,
103'h1a3e18ecac641f870801f0c765,
103'h168b71261e69a5acd200000000,
103'h20d44d1fb8a7be998000000000,
103'h2afc07194f332fbf9e00000000,
103'h3d419d1b31077cdf5600000000,
103'h3ceb52a41a0383f8a400000000,
103'h1afeadd9d6452113d4001fd5bb,
103'h30b9c7a9143073b7ee00000000,
103'h16a81137ef2f2191c600000000,
103'h2a9dd7a620e8e93ada00000000,
103'h1a97220cf690fa72c804b91067,
103'h20d58d87a02ed218e800000000,
103'h3a446cba3ac5f425de00000000,
103'h02e26d7e9a9b81ad807136bf4d,
103'h2c69577dd4dfee67ba00000000,
103'h0a813befd8c25be656000813be,
103'h0ac7f27ac42bb3642a0000031f,
103'h06d49d2b8eacef540200000000,
103'h1d7cc989da74e1cec600000000,
103'h0704e44fe1497efa5600000001,
103'h0b4f5afc3cc6488430000000a7,
103'h10c5850cc2cb2cd410fd2c1c59,
103'h26e89e714d1a87d04c00000000,
103'h168099a49ee00cdd0e00000000,
103'h266213d244c8ab4e5c00000000,
103'h3309d6841d4944f2fb00000000,
103'h027cc60a02ab58c53e80000000,
103'h1f0a3d6036b52f495a00000000,
103'h1977c1937931f5535e00000000,
103'h16adf115173c32b39400000000,
103'h332d6589aeb3f4470d00000000,
103'h105832c38561e55c227b26b3b1,
103'h24382f46b68f4ae5d000000000,
103'h304a211d46e77da95400000000,
103'h129845a76b1facf00c00000000,
103'h229a5e789a69ce0d5200000000,
103'h36fe5ca5ed0213b4be00000000,
103'h02f1a5b90e9c722d582dc87000,
103'h16cc6c75869aced34600000000,
103'h14c6e022088c748c5400000000,
103'h2c2b21dbde58e101da00000000,
103'h3291774a731fc123e500000000,
103'h08943ee6604ae2ffc26f6e0cd1,
103'h2231d55592dc5a4a3600000000,
103'h065be0511b7099309600000001,
103'h0adecc4e7ea26e8628000006f6,
103'h0081796fc4fe4ed744bfe42384,
103'h166f0990cedd1b25c200000000,
103'h3e38f3fc0e5e94958600000000,
103'h02737797e4cd9e2656de5f9000,
103'h055069b9e40692226400000001,
103'h0c2baab3277a09ba4abdd5ddb7,
103'h22e406d22cca73742e00000000,
103'h06faf786b8f61e275400000000,
103'h10df86619ada24f98002b0b40d,
103'h3ecaa75ee0d51c803800000000,
103'h152fd21672b4a2e1d200000000,
103'h145f7042317f4a40b400000000,
103'h0e852c9544af1c572642860a82,
103'h20850de1da0e8c995600000000,
103'h155a0baea893b92e9c00000000,
103'h3ae3ac5d4918c7107700000000,
103'h12ec974c9f72d2bf1e00000000,
103'h2ea49e9318567f1c6600000000,
103'h246b3272ea4316690400000000,
103'h02c57f8158e7b4fc1ee0560000,
103'h283893a03c52e76f0800000000,
103'h2e1e7a7e3f1866f06200000000,
103'h0d5ae078a850fa909ead7d7c5f,
103'h14da5cdc176f750ede00000000,
103'h37418e3ba2ca55878600000000,
103'h16fba70a36a4b2639c00000000,
103'h34ce26c92ee6409f3e00000000,
103'h3af1a118c4e1e7a97500000000,
103'h1684907738b00e72a200000000,
103'h14e1d55d32a1af8b6600000000,
103'h08e3cca6c82640029e62c6522b,
103'h2ccc048f9c08155fd000000000,
103'h12962421e4ebe2069800000000,
103'h32105226d0b7e6963500000000,
103'h032c2fb7254e0ab81afb724000,
103'h1d6e4d4a165e5cdeea00000000,
103'h10b8803cd88a8c960e16f9d365,
103'h2aee953634f8d9e02400000000,
103'h16dc90c5c6b15a1cfe00000000,
103'h2418970d709fef533200000000,
103'h0ab2fa34067c8018f800000005,
103'h08d7e9f0ac9517266a217f6b63,
103'h3af5b38d7648115a7100000000,
103'h34c4d7473e1ffb4b1c00000000,
103'h1e33ea543815aed89200000000,
103'h0e1f7d7a2cda861fd00d020d00,
103'h2ca027c68b0e70740a00000000,
103'h3f68e36d5a2dedee3700000000,
103'h11519a5f46ce15b4c241c25542,
103'h1a500029c536f9221c0000a000,
103'h1028ec141488938162d02c4959,
103'h121048726ed893ab2600000000,
103'h2f2592bf01017fbf3c00000000,
103'h1008f2c05211c831aafb954754,
103'h39234be3c2375af0ab00000000,
103'h34c6388893404db0fe00000000,
103'h1e41b8d88b639994c000000000,
103'h0abeb8e7be29d21d52002fae39,
103'h094d81289f6b8af5de1305eea0,
103'h0913a45a282a43dd9c9cf3c3da,
103'h1b1a153cb077c5063afffffffc,
103'h38841fb3f88b69606300000000,
103'h1617fc4892a57e9d1200000000,
103'h111763d30c299e510a76e2c101,
103'h35410f3b23419a999e00000000,
103'h06e27fa97358fe6caa00000001,
103'h120f5978269a0da7cc00000000,
103'h30e1b1e3ee7c8d513e00000000,
103'h1adda8a0c08be6c96600000dda,
103'h271b39f7316d98ad5400000000,
103'h24b1c9ba4b4b414e1400000000,
103'h0ae2672531667b45441c4ce4a6,
103'h1e8f91e1551844ff8e00000000,
103'h32c8a366e0faac24bf00000000,
103'h366f4d99be8a3e061200000000,
103'h0561391ab252e16cf200000001,
103'h02b99fe0e8c22f06b2e8000000,
103'h172a4ba6af2368216400000000,
103'h0895a39130dd08024c2455c9be,
103'h3a8b3981c60753a8fb00000000,
103'h1ed3b0df509cf73a2c00000000,
103'h2cde57438a2830bbf200000000,
103'h270c65c92afbe19b4200000000,
103'h13177c5116da38dece00000000,
103'h0629e681fce69ea7f800000001,
103'h08d947ed10fe1af90e13ae8a0f,
103'h16b0da141628017b0a00000000,
103'h0e844dd65e0149681a0024a00d,
103'h1d31fa7776b2237c3000000000,
103'h28c645c0853671529000000000,
103'h0358ac02a3686bca0662b00a88,
103'h351313bfca2eb18a8a00000000,
103'h04cec4e50c875d8d2c00000000,
103'h0a3c9986809a714cf600000003,
103'h14e0df7a856936320400000000,
103'h02ed91388ea5cfb884db22711c,
103'h3928f4812486af330b00000000,
103'h3cebb556e674406b9800000000,
103'h0248e7799e9d34ecbcc0000000,
103'h0d0f4fce5c88ea43a2c7f7e7ff,
103'h257b87db9ed1d1bd4200000000,
103'h236e6f1beae1218b9e00000000,
103'h04d596c7cf5ca9673c00000000,
103'h06d9f36070cb18832600000000,
103'h25673a3cb6a0af4af400000000,
103'h20c652d63d7aa2ab6600000000,
103'h07068cfb62e1dce81c00000000,
103'h3ca37087c2a82fbe5900000000,
103'h230b6c974aaebcb9ba00000000,
103'h3f1417f1c7522d417e00000000,
103'h169765f7a95d99d8c800000000,
103'h12fc90e5a771b1ca8e00000000,
103'h1009eb91fd0917c2368069e7e3,
103'h18c602f80f05a8a7dc00000000,
103'h26d4479f9e0f9439d800000000,
103'h1c40261ff6d59731e800000000,
103'h381db66adca9ded18700000000,
103'h10045e77f8ea04f17e8d2cc33d,
103'h38f0af2cf007bb5c5a00000000,
103'h00ec941bc30c19d454fc56f80b,
103'h3ebe103c7afcc9014400000000,
103'h18396b2ebae95d1d0600000000,
103'h2c9ecb1278a76d598200000000,
103'h330be65292e0d8883d00000000,
103'h38851b66ff7fa39ab600000000,
103'h3afb197cb08b89ed4900000000,
103'h395a74af6a10a5544700000000,
103'h2e613d3ba50bbed0f800000000,
103'h3648de501d6633806200000000,
103'h3cb022ff4ac770bc0700000000,
103'h34a2f19bc1104f0c2400000000,
103'h16a6658c7ec0720b6e00000000,
103'h1eb5984e336363a73000000000,
103'h032afe904b09c933ae12800000,
103'h3167d58e68bf6181e000000000,
103'h20b4fb98aaea60122a00000000,
103'h0ec293ae5a5235a0922108d009,
103'h31338f6b3c0731393c00000000,
103'h1aae545bcac9c4e798000572a2,
103'h2ee87ace3afd5452d400000000,
103'h2b0d0152d6aba8ae9e00000000,
103'h0283bd780494237cdad7804000,
103'h1601aad66ea124cfb000000000,
103'h37495d1c7324e247b400000000,
103'h108e63b548268d1e2233eb4b93,
103'h007f12fcbe6fea3a94777e9ba9,
103'h3403e5c10efe4defde00000000,
103'h1629dd550e7d60ec9c00000000,
103'h2c74b730c28146adac00000000,
103'h0ae61e2a9aab2402ba00000003,
103'h26c76f5f071fdb337e00000000,
103'h12a70e835105f95e1800000000,
103'h0e040e9436cd68bd1e02044a0b,
103'h0ce25552cb7477406efb3ba977,
103'h256bc014187885d4a400000000,
103'h03150608e45adb276e39000000,
103'h30c4455bc8c69b3b8600000000,
103'h1540ed6bcadba1446a00000000,
103'h05320cbc3a9fe6a03200000001,
103'h0a9bb1e14ee0d40bfc00000001,
103'h3660322dd212e0c83600000000,
103'h28eb4db5deae92a98600000000,
103'h27520a82540ec4d75800000000,
103'h1c58adeefcfa128d3600000000,
103'h22402567a24c1d0f8a00000000,
103'h3d3a7da880a4cafe8800000000,
103'h32e36892e2e4f0662b00000000,
103'h3e9b18549e1f6e0eab00000000,
103'h074cdaa39302d6a18e00000000,
103'h314aba02109deef62c00000000,
103'h1ced645f16eac999be00000000,
103'h2a74ff224635839bce00000000,
103'h161c07f42222e7fae400000000,
103'h16c5e7678c97e71d2c00000000,
103'h250db5d124b3ef114e00000000,
103'h0b404dd47b79d678dc0002809b,
103'h36a869739e878c4a0000000000,
103'h04336d0da8c7da1e7a00000001,
103'h205657c4de7043921800000000,
103'h212d318d64a3b09fc200000000,
103'h1a7de1cec4fa0864a000003ef0,
103'h35561e5a262739f20400000000,
103'h36f6350400a51bc0ca00000000,
103'h16068f3ff4fb3a1af000000000,
103'h1cba9a1baaf16f1ef000000000,
103'h2768ad5c02f7fe5ee600000000,
103'h173dfa8e5eb2987a9000000000,
103'h06b86381841b45d69200000000,
103'h2d2e068f9a594064f000000000,
103'h3e9518bca011a3e67500000000,
103'h10f429488e3faa760e5a3f6940,
103'h0305d24f0cd4c332b086000000,
103'h3632c12c1cc8ec7b3e00000000,
103'h06b8f06e1ecebeca4a00000001,
103'h3750c39696017ff66600000000,
103'h352841351cba70648600000000,
103'h3ed48206530b33fb1c00000000,
103'h2549af52c73375303800000000,
103'h2a8d9b698507f7368a00000000,
103'h06d30776a951a6895000000001,
103'h3ed2e3e854df41f2d400000000,
103'h08ddf4551ab249697c37de9e33,
103'h191c79f21a852d51d000000000,
103'h2c62f6c5a36321a6ec00000000,
103'h2afb1a227d7f9b990600000000,
103'h3a727f7228e2925ea800000000,
103'h269c2e2b52ddac812400000000,
103'h2d4b0a364f502bf34e00000000,
103'h165d07e834ec5a1ea000000000,
103'h3aeea13322376454ef00000000,
103'h0962ccdcb8946c3d24fb5070ce,
103'h2ab4a50772830d704600000000,
103'h1956a9257ce5da4cfe00000000,
103'h3ce50762269a7f547000000000,
103'h02aac9f3bef12879ec77c00000,
103'h0104f8c27cd62fdc12ed944f47,
103'h32e235017e80f9cfd300000000,
103'h1ea54b8d8085f2924e00000000,
103'h3302e16df2682793cd00000000,
103'h04519fc8500d73214c00000000,
103'h12768dfec210548f3e00000000,
103'h1e1c76050761f4579000000000,
103'h2c48509d98d882565200000000,
103'h2adc52c9f8f4f85b5a00000000,
103'h3b7dc817a43d48f8f200000000,
103'h0e2f91f48e199bc2ea04c8e045,
103'h294350290a9763da8e00000000,
103'h1b2f90b3d8c6f5cf1effff2f90,
103'h0710c99a010a45f82800000000,
103'h142f4b791b39d6ac0000000000,
103'h3267691b214aa0460100000000,
103'h1b36ea97b679ebbf1afffcdbaa,
103'h1acd61e368e154da3c00000001,
103'h1b6e1f2745183f71f2ffffffdb,
103'h3648b3171ee5a1555a00000000,
103'h336de74cfa53c07c9f00000000,
103'h250d0741f09c7393be00000000,
103'h3e8d7c11230a5ae0b800000000,
103'h1f26305247176222a800000000,
103'h1ca485e8c4a4de33ca00000000,
103'h14769bfbe2cb0e861000000000,
103'h3ce525a2be6f946ed400000000,
103'h065e0a2a52e6306ab800000001,
103'h16ee50d48ecb560d7600000000,
103'h2a2375b295296037ca00000000,
103'h2223a916aa17b10c5800000000,
103'h1a9370e9973b26beee00000093,
103'h24e96927385ecfd59800000000,
103'h3c0ab77252f240bf2f00000000,
103'h2a5565f536dba9e66800000000,
103'h04b7c58474e66158ba00000001,
103'h32554bd29f3bc74df300000000,
103'h1a51a1f662f38cd2660000051a,
103'h174038d95648d8a50400000000,
103'h080a79a2b09a7a9b6848019cec,
103'h2ebb1bc4c6dab374be00000000,
103'h32a78534cee52d176f00000000,
103'h1a877b773ca048dc3600000008,
103'h18b04a5eb047ce110400000000,
103'h087393e18acf4988425e6d34e4,
103'h3f1190d9257f93e6f200000000,
103'h0294bae82cf327c87c80000000,
103'h04b82dd36a04b8a1a000000000,
103'h36236ecfac997389cc00000000,
103'h355df9543251a15d3600000000,
103'h141817bfa975102ce400000000,
103'h22c55df39cd309811600000000,
103'h19775cc932eb2140be00000000,
103'h3cc2cf2894b07f345c00000000,
103'h125fe2e52d27dbfd8e00000000,
103'h137206ceaaeaab262200000000,
103'h2e5734393c4a8e0b4e00000000,
103'h3c2782e48ebc94d9f900000000,
103'h1ea850c43d13c9133600000000,
103'h2c50faa1783b4bf7c400000000,
103'h26e44fa4d6e39cbc0200000000,
103'h1cc232b38434975d7a00000000,
103'h215caa9c2b18e7025200000000,
103'h230aeb9806db19b5d600000000,
103'h1ef4788ba737c4520000000000,
103'h30c1a23b4b42afea0600000000,
103'h06c3634868372875ac00000000,
103'h06de0b57d8f8cab0f600000001,
103'h0cd3cd1d1ebc2df95e7ff6feaf,
103'h39015334649a39513700000000,
103'h31718935b06e066e5400000000,
103'h0e18e7aca86f59a2b80420d054,
103'h06b910d498e0e2d86800000001,
103'h1b1567f5e8f9ca8512ffc559fd,
103'h150bf8686eb2db59aa00000000,
103'h3c708f4948c8434f9300000000,
103'h0e447fccdcd43bb800221dc400,
103'h3af95328db44cb014b00000000,
103'h0ca7f109e8894ace2657fde7f7,
103'h0e096a44a2829df70000042200,
103'h193326cef12a8f00ea00000000,
103'h3f311f113e33f9458d00000000,
103'h0173e254d66720147ced8134a9,
103'h2a3ff06694983f25ba00000000,
103'h368e9c6f540c217a9000000000,
103'h3407d778ff4c11e12600000000,
103'h2eb50bc836daae507a00000000,
103'h00c9602beae285c97ad5f2fab2,
103'h2675f3b558979191b000000000,
103'h202ea8b95960f1bd9a00000000,
103'h1a336f9e7ed6e572f20000000c,
103'h0b12e4d421058e2c4c0225c9a8,
103'h24d4dfd33a38fdcaca00000000,
103'h192e6c64064be29eea00000000,
103'h24e8eab26b20c2722600000000,
103'h2e7a4e73c34f2ed62c00000000,
103'h1a114061663819889600011406,
103'h00e13019d6b267fc5ac9cc0b18,
103'h2cfd027130c3a85dc000000000,
103'h0339973ab0a4d877965ceac000,
103'h1cc55ada5ca1dae8c600000000,
103'h1e8938029edb72237600000000,
103'h34ff7d273ca0ccfdd200000000,
103'h3d396aa99b2a05007200000000,
103'h321830a38f298227af00000000,
103'h0698d1864b62ecd14800000001,
103'h38f4e48c7e7b1d74d600000000,
103'h26f1c4908513eefb2200000000,
103'h2f18a994fd08d387a000000000,
103'h056910c122fa98182400000001,
103'h271c64be911341ad2000000000,
103'h064ad630d57c526e4200000001,
103'h2a8d369e3c98b72cd200000000,
103'h0ad86a9342e38d5da600000d86,
103'h0d1e36a06e70c3fbe2bf7bfdf7,
103'h1e77445ab9492e8f2600000000,
103'h074ca4834767652f9400000001,
103'h28babbd8a4dea98a4c00000000,
103'h0e0c608baa2b4e0d92042004c1,
103'h22cec93a94e609e63800000000,
103'h30da6078a2f26a71e200000000,
103'h034d5ce646c133ac7618000000,
103'h3a9f02de369b94251b00000000,
103'h1e1bf6e3b8e8f10b6000000000,
103'h157ef4cf7487f3e99600000000,
103'h2ed45d2d12a3eacd4e00000000,
103'h0eeaf9372622df9cc2116c8a01,
103'h249d296656f73cc9d400000000,
103'h34384aa0e4e23600fc00000000,
103'h375b5fc50b7f5f675200000000,
103'h0d225fb67eb7aa0836dbffdf3f,
103'h080c3f44b41309cd400f9b44fa,
103'h1aed5b9cc0356983be00000000,
103'h10b0adf5c941a8c874b78296aa,
103'h12f35fb6222f04653400000000,
103'h10edbb7eb4dfb25afe070491db,
103'h04fb211486d312112000000000,
103'h3a3df02e16c0cd8fd400000000,
103'h38c268101cbbeea45a00000000,
103'h1975e45756f9ded27200000000,
103'h2f0912f98ebc46e28e00000000,
103'h086f53ace7322b39e4aebc4a81,
103'h3a9661f0153b3e337300000000,
103'h09795ed79eaa91e058e9e79be3,
103'h2c563a919940f3d06e00000000,
103'h1eef5d2e22ba52a80c00000000,
103'h38baab048e108d39a400000000,
103'h26c1370e6effea67c600000000,
103'h337254f8a6ba956c5700000000,
103'h176466b34d7bcc7ac400000000,
103'h1f10cb15feee21736a00000000,
103'h34cdbcb255528826b600000000,
103'h388a98b67363533cb400000000,
103'h22020a26e6310fef0800000000,
103'h18f548121ebba8a57c00000000,
103'h0cd6a770c0bdb2cc627fdbfe71,
103'h140a8ef618b2fade8200000000,
103'h10a1c9b82489a24f420c13b471,
103'h356a14693a9431455c00000000,
103'h36ee07bfca35fafd8000000000,
103'h382fade2bea00f66bb00000000,
103'h14244ee4348e17268600000000,
103'h16a29234eebdc5094400000000,
103'h10b506cb02e213ed7ae9796ec4,
103'h16fd765e9884a6226800000000,
103'h1ce5f558ea39aced6a00000000,
103'h165c8b79c137234c0400000000,
103'h3e90e6a3dd1d18a4ee00000000,
103'h28a755bb7279a41eae00000000,
103'h2c426af5710a8ac28c00000000,
103'h1b172d1cdab1e07dfeffffffff,
103'h0a23129046f44b737000000011,
103'h174c10a8a30b78904a00000000,
103'h14eeb2dfac2e8b209000000000,
103'h049bdfd9427a9bc93200000000,
103'h0efaed50d6694ea8de3426006b,
103'h214e463bdc052e822000000000,
103'h12ad17b72b001bd2f800000000,
103'h323a74530b4e620ed500000000,
103'h13426cb81efb79c5fe00000000,
103'h0ab3b3c61135ee190a02cecf18,
103'h1e2a295623785ad12800000000,
103'h1ea0bab92f2c0e973800000000,
103'h2865ae2b0c5637ed5a00000000,
103'h10261b62eaf6f2a68897945e31,
103'h081c76b3d35ca0d196a06b3122,
103'h228b2cd5e282bc348000000000,
103'h2c25f18f2a9f32e85400000000,
103'h0316ee35ce2a5fbe3638000000,
103'h02fedd82fb50514d6282fa0000,
103'h17436da1bd673f833000000000,
103'h0e0ab9f4ff661d062a010c8215,
103'h3171393096a98aa7e600000000,
103'h2102182a64b4449ce400000000,
103'h0ae3487194257dcd7a00000003,
103'h312bb83bf42795f7de00000000,
103'h14da450c7e0ade697200000000,
103'h11325c84ee3696a5667de2efc4,
103'h2e3eb89a4210dbb1e400000000,
103'h2270927d12433836d200000000,
103'h08ca0257c281f0d11625f9436a,
103'h2f2e509be4f2834e2800000000,
103'h00c935856cbc85a5eac2dd95ab,
103'h1674f620daead641ce00000000,
103'h0163eef31cb40bc73c0bfd5d2c,
103'h2ad4d896722901e81600000000,
103'h3a384587f28cf0db3200000000,
103'h3758381f5f61c971a600000000,
103'h0d6300f8989a0ef998fd877ccc,
103'h0121d5990ef24718f60a0e5902,
103'h2609ac219a5548118e00000000,
103'h3e7e73855a771daa9d00000000,
103'h3655045ac080c9cc3800000000,
103'h04c5a429c0ff3d519200000001,
103'h23288b11b75441ac5400000000,
103'h1ae0ba0b3b19e5d614001c1741,
103'h2c1006af5d4270e7ca00000000,
103'h00c01d1fb6232af30471a4095d,
103'h156f70e1a53331a26200000000,
103'h1e73064fe4f34ec21800000000,
103'h249081943a62bfa3bc00000000,
103'h06f06dc058d5c5f3a200000000,
103'h1e7384df7d664787dc00000000,
103'h1c29cda10256b5483400000000,
103'h3ed36524a2ca3a27b300000000,
103'h1adfbc4bfef407c8b40000001b,
103'h0ec1d966fcc76ced5660a4322a,
103'h010a3e09d6a7293954d8b3a195,
103'h36a957f4e46902a05000000000,
103'h0d12ac07a67340aa26b9f657d3,
103'h237007e31d1c989f0c00000000,
103'h3294d0abe92f44a6b300000000,
103'h1a60c2ae0a9f4c89ce0060c2ae,
103'h2695b7507e341d35b600000000,
103'h193dec9d1894dfe3c200000000,
103'h2702ba88bf2a97344000000000,
103'h1cf6cd1b176883d15800000000,
103'h1e8a2c373d6b3e5a1600000000,
103'h1e51a88919620b752c00000000,
103'h36ae04beb8ec37ac6800000000,
103'h0c34f828963de035801efc1ecb,
103'h39246f63ceebe4f43900000000,
103'h207f24f91b20dd1cd000000000,
103'h233be60395454c809e00000000,
103'h1ae4deba74c47179b800000007,
103'h2acbb7a6d600577d4c00000000,
103'h089e758772e53637c23da1d858,
103'h02921084dcb0edde988426e000,
103'h0ecaf802e64f63660a25300101,
103'h10c850faa8e173eae8f36e87e0,
103'h2ac6016fb6ac6bedce00000000,
103'h34a8e81c8974bce87600000000,
103'h1d3cbca7f23abe582c00000000,
103'h2a1ff49966e3a674b400000000,
103'h20e4a075c420631ca600000000,
103'h0e55b83fef4057b60e20081b07,
103'h033b8cf29124f82bd28cf29000,
103'h2b5c1ffd5e7ab06bc000000000,
103'h3860597ce0b63d5e5100000000,
103'h0a84f6190a125d5bae00000084,
103'h0ae9ea6b4372b6d8900074f535,
103'h1c73d6e94cf7acf19a00000000,
103'h0b7873d318e1975cde00017873,
103'h1b334e1b34556e462afffffccd,
103'h360085befecde2194200000000,
103'h1540743b5a0130347600000000,
103'h3f780fa95101b5f37700000000,
103'h0291427425422a2ed0a13a1200,
103'h38ffe38522ba39d82000000000,
103'h2e3c66af654b7c4c4400000000,
103'h3f7a1a0e1e4b5fd16700000000,
103'h1eb983604c87c680cc00000000,
103'h233b16e14d01e08eea00000000,
103'h0a76e43a6abb63ef3600000007,
103'h16fe2ddfcef67ad08200000000,
103'h00d0d756996d5f0aee1f1b30c3,
103'h372b474e2f6b8ceabc00000000,
103'h3a8797d4af3c64415500000000,
103'h289f4c4a6567ab8f8200000000,
103'h24ad7b909eef43643000000000,
103'h382909e1c68e8fae9500000000,
103'h3a10251dab3c0b3f3500000000,
103'h2a33a49ae2651520fa00000000,
103'h3ebecfa79d753a3ea600000000,
103'h32393e1886a8ded98900000000,
103'h2f423c380767ae812600000000,
103'h14874596b8a0ec99ac00000000,
103'h1c31641666e328d1b200000000,
103'h0250bcd4bb6a6e686c97400000,
103'h3118f46c989bd27ed200000000,
103'h2248da859aec8f538e00000000,
103'h0e19ad384b0583c02600c08001,
103'h22cda8bcae4e5e45c000000000,
103'h30ec12a97d680b7e0c00000000,
103'h16a64f151f35b43aba00000000,
103'h164d1ad44e21c6e43600000000,
103'h22f96a53a4c815f95600000000,
103'h1cf41818bc1530cda400000000,
103'h1456d15bdf0e9b214a00000000,
103'h2aef3ed9bd02b33a0600000000,
103'h0ea9733bd0598495e4048008e0,
103'h192bbd973a48c36fa000000000,
103'h1ec338c048f236ab7000000000,
103'h05694f0aa21df442aa00000001,
103'h2412188f00e12d02f400000000,
103'h161466a9454a7c0d9600000000,
103'h015f78332a5c949c96de0667e0,
103'h349cc0688170fb45dc00000000,
103'h0af7fce080d07379060f7fce08,
103'h2334665b776d33e18600000000,
103'h3ebb4be4006530c20700000000,
103'h049ec6092299971d7c00000000,
103'h0af33b742154e3017e00000000,
103'h1018245824f3a90aa0923da6c2,
103'h0eaa411daee6e47ec251200e41,
103'h0ca18ea540ff08d6e67fc77bf3,
103'h2d32734a4ea949f49600000000,
103'h2f183af0db4ad899d600000000,
103'h16f1aba2077d4be42400000000,
103'h2cb200d1f69586d4fe00000000,
103'h03715ed8cc87327704e2bdb198,
103'h26da06d438393348fa00000000,
103'h248d87697aaa9221c600000000,
103'h28be53e2e08498f5fe00000000,
103'h2484a7314412205f7800000000,
103'h2ad22cf6acd074425800000000,
103'h2a58e60510551b739c00000000,
103'h228a31353d27486a4a00000000,
103'h3d40155b66802e6f5a00000000,
103'h180819e1080a5fa49600000000,
103'h22a092a9044a74fffc00000000,
103'h3e8e26e49f528ee10600000000,
103'h14a3038a80f3218a0a00000000,
103'h12380e9fbe81486ea800000000,
103'h18d7795995244bf92a00000000,
103'h22c15913665c5a98e800000000,
103'h0cfdc7ae3e33d3f27c7febff3f,
103'h362d57d320f52d05e200000000,
103'h1ede3066acf2f4b42000000000,
103'h1cb354f363204c874200000000,
103'h3ee4d41902fe7cedee00000000,
103'h214a27311eb1d1e15200000000,
103'h22a4a74f1c96a5fa5400000000,
103'h10f21c213ce0cd2b7208a77ae5,
103'h225fdd7a9e85747a8e00000000,
103'h36cc1bc1f177909bcc00000000,
103'h28ea2bea92d76e166a00000000,
103'h389ee20d8aa389d85b00000000,
103'h0434655bf28db5c2ee00000001,
103'h2e4f5d24eb2c97d07800000000,
103'h0ae1e589ae60fd2c6a00000387,
103'h394bdc04deb05a515700000000,
103'h31595c5868923fdb0400000000,
103'h1af4926ee0de1bdfe200003d24,
103'h30bc6055d03778384a00000000,
103'h36e52b692a2c0aa72a00000000,
103'h18be50cddce86afcfa00000000,
103'h2529b60d92cd96662600000000,
103'h0e73372d2a8be7340201939201,
103'h0af430850eb59d4194001e8610,
103'h30a134841e28d46ebe00000000,
103'h3336a380291d04f3cf00000000,
103'h0699a8e258be3977ec00000001,
103'h048895788af4dcf81400000001,
103'h132d1f50508e85da6c00000000,
103'h3efa7d96d5171b52f600000000,
103'h12e4e0d129443aa34600000000,
103'h3e8d7d83663eb83a1b00000000,
103'h352af72dba23990b4200000000,
103'h3a56f6b278b1168eaa00000000,
103'h169a118a2edc0dbc6400000000,
103'h182167052833046edc00000000,
103'h02e774ba3ecd15f90a774ba3e0,
103'h26d11b7a98ee7cfe3400000000,
103'h046bd8c99ad5f1b87200000001,
103'h0ee2a3d502a70d330a51008881,
103'h028c734f4712e5fca63d180000,
103'h360358c294f589d1a800000000,
103'h0168bb341881fd20eef55c2a83,
103'h26a40f5e0e8555e38200000000,
103'h0e8670bb0eee11179a43080985,
103'h3d7bb814b6922075a800000000,
103'h0066894005189130b8bf8d385e,
103'h1ad3578c429449456e000000d3,
103'h04c57bbc02fad2857200000001,
103'h3ca5b1035cce2a11b500000000,
103'h2a1806c06093a5cdb600000000,
103'h1ca2edae1d3956d11400000000,
103'h12c21de146515d917400000000,
103'h08dc2099e4f44b3f921435d33b,
103'h1cc44d6436b66920d800000000,
103'h12401ffc3e9289babc00000000,
103'h24f549655c56d71ef200000000,
103'h3cfbd05fee96f71b3200000000,
103'h3af6a29a128c40808f00000000,
103'h2ca7ddf50e8810e07c00000000,
103'h1eeba30ac97eb37a8e00000000,
103'h2c863f3f7626916f9c00000000,
103'h28b7d28f5512347a6600000000,
103'h3775a65fc29873b9dc00000000,
103'h14bb8b10aa5046493000000000,
103'h3a80233c22c5eca8f200000000,
103'h176b4cd7368177b99e00000000,
103'h0768aaecb1019af5c000000000,
103'h3afe7cbc076ce7ccf700000000,
103'h18e494d48cd592b9a600000000,
103'h1890999606d40f75ac00000000,
103'h0ebe16111eb8a44a385c02000c,
103'h34ed2d81f7493de04000000000,
103'h20892cbfc40753f15e00000000,
103'h18fabeb738f481735600000000,
103'h18406024587dae331a00000000,
103'h393ea5dbb3786cea5500000000,
103'h0e8629734ab8cd0eac40048104,
103'h28d500fc42f772ea5e00000000,
103'h3c1859f8917d9c5dab00000000,
103'h2ad96127fa529d59ec00000000,
103'h0812d541b76af7527ebc1109e4,
103'h3205166a2144587a7900000000,
103'h20eeca7cea572dbc2e00000000,
103'h1e561aed5d5c44265000000000,
103'h161008b7bd4b0ea33a00000000,
103'h0434edd49aa129909600000001,
103'h149e2b6bf0b132485400000000,
103'h0f5e96bf76e6201cee23000e33,
103'h267b46394a844b88e000000000,
103'h3ae304565ae2e2485700000000,
103'h28ebec04005e2881a000000000,
103'h08a605f9fa412cd7fa73949700,
103'h1e46400ce22d18dbfa00000000,
103'h016ac5a8acd31ed5f41ef23f50,
103'h3a722d8ccb195ee2d900000000,
103'h36d7bdf28a84248b8400000000,
103'h2b7e7b3046f652184e00000000,
103'h03525149fcce100ada149fc000,
103'h06f94639a74c8b3b2000000001,
103'h16b99a0c2a9edc851c00000000,
103'h30fe126a309822bec200000000,
103'h1038dce08651bccaecf3900acd,
103'h2c41b761b74fcf351e00000000,
103'h2e971d1e0688ac15a400000000,
103'h1c8b5f5f72ca63775c00000000,
103'h3b17c45fa26180956200000000,
103'h1ef5e62abeecdff4d600000000,
103'h3b23d72af904a4547900000000,
103'h1eda7440d6fa8a7f3600000000,
103'h355b74ce131e61aa2e00000000,
103'h2d3df5f0b0f8d5eb0400000000,
103'h230d570824544ab91600000000,
103'h10e15c74109240a9c6278de525,
103'h14afec5f329f97b1ea00000000,
103'h2c9cddf48280f425fa00000000,
103'h3282a574d630e0852d00000000,
103'h1ebcb7ae42cdbe79ae00000000,
103'h18890a91775063ee8600000000,
103'h06f4f526940d1b9cc800000000,
103'h34e1d3e1ac96262e3e00000000,
103'h3aff9321f28b1b54d300000000,
103'h04eb10dbe96cef368000000000,
103'h0226f284626c82587262000000,
103'h166fefc9a65793345a00000000,
103'h174f133d2b7e85b8be00000000,
103'h08b9520580ee7582642b93c3f2,
103'h24908004563d88bf8e00000000,
103'h22d4305b9ef6dac50e00000000,
103'h066f73e742875ac96400000001,
103'h16893d2ba55b8b250400000000,
103'h24917bf26ccaff0c4600000000,
103'h0ad74378c3543c37ec000001ae,
103'h0e13e5c426e5b82a5800d00000,
103'h14d7e2d8f0bcfba31a00000000,
103'h00f76b12bed0e16740e4263cff,
103'h18e1f258d4a8c4403200000000,
103'h3220b5d6d4a02f52f100000000,
103'h3545317f2e8221abc400000000,
103'h2626a8caa0a2d7829a00000000,
103'h16d9017d54e80901c800000000,
103'h1c341e703a0eb1cc6800000000,
103'h372f6ab612e7b349be00000000,
103'h3eacd8a7ae1bd1b9f900000000,
103'h26cd1e1be44b3c700a00000000,
103'h24d56c91e2f81517b800000000,
103'h1eec6cd448c533339c00000000,
103'h28eb20606e9a9fc57e00000000,
103'h2305a5a68c870c99c800000000,
103'h3e6b675cb5722cfa3600000000,
103'h3ec93e2a9777d2a0c200000000,
103'h06ec482c16e339fd7600000000,
103'h3ca9f1f314ac78280f00000000,
103'h3eeea853da98c0542500000000,
103'h34a58baed742b2473800000000,
103'h02d441aa95315a9b1241aa9400,
103'h26e631a3c8d6e649e800000000,
103'h1ea499c50cab27f47c00000000,
103'h30fbc23a729159984400000000,
103'h18959cf71235f35d5000000000,
103'h1460d24ec331b597c400000000,
103'h1b02edf05cc7528ed6fff02edf,
103'h2a503186702824dd9800000000,
103'h2e2eceb4ca2b12cdf400000000,
103'h05435f40777b44546600000001,
103'h1e89a563e4aa13093000000000,
103'h12973e162aed7249a600000000,
103'h38ccfba6097717ad8c00000000,
103'h2a2dcc03db0e55c3b600000000,
103'h1109e0b614db5169be1747a62b,
103'h1c9008717e091d6d9800000000,
103'h1203a2768e12fe23ac00000000,
103'h10ee54292ca306952a25a6ca01,
103'h2ae75b9f7ea6a90bba00000000,
103'h16bbb47f9094fd34e600000000,
103'h02992acd3a7c58d4649a740000,
103'h3c899f3e90380d53f400000000,
103'h221d1a4512d138212e00000000,
103'h06573e574f5ad75fc000000001,
103'h3c265f9e7077f1a4d300000000,
103'h2b71d9b9f8cf2ffc2200000000,
103'h2af5612974f58f9a9200000000,
103'h3e4a20ba1e6769548a00000000,
103'h20f9b7aa8a5cca7dfe00000000,
103'h3321403fc8a6eb381f00000000,
103'h3f17f8d128a0a2e2a900000000,
103'h3c0440fd1ac1e3227100000000,
103'h1a57f27d98d9dbf3980002bf93,
103'h03086e7c16de1cf0b216000000,
103'h325fd5b2b1360f6e4d00000000,
103'h0b57dfcbf53e7dea62000055f7,
103'h3e11cd07a69e539d1200000000,
103'h0aa59636f2f63369060a59636f,
103'h2d177c56f1080070ae00000000,
103'h3ebf71e53aad96a7a100000000,
103'h06a5e55de6c512fe9000000001,
103'h342aac73a48484e3ca00000000,
103'h14a5a6f26b2a6a41b000000000,
103'h2428a1e1de5516b55400000000,
103'h2e593378f2fabda7c000000000,
103'h1e4ed80e96235f899e00000000,
103'h32c90188057c93029300000000,
103'h326d954322cb6b112900000000,
103'h13673fb396946c992e00000000,
103'h245ba7cbc80201dc5000000000,
103'h0c736f6d9a69418fe63db7f7ff,
103'h3a07ca11fec4e95bb000000000,
103'h0d678fc78c3858c94abfefe7e7,
103'h325bc216474022db4b00000000,
103'h2251f64152a7b2a2d600000000,
103'h2eb16bfc460374b91c00000000,
103'h38d5cb12e9556afa7000000000,
103'h0e3282f2d706d6f6b60141794b,
103'h2acf5dae0edca2099e00000000,
103'h1a13eb0c1d0f24fc7600000001,
103'h115bed2348de82aa843eb53c62,
103'h30f95a34e2f26db6a200000000,
103'h269d9e3d354e5ad9ea00000000,
103'h2b1e844f2447b50ecc00000000,
103'h0cae8f5d8ae5534c0077efaec5,
103'h361d1d167403d79b2400000000,
103'h057e188602b266f8ae00000001,
103'h042d6ecf78cf840f2400000001,
103'h2a247a27bd4d9c952600000000,
103'h1900d8cc027b0b649e00000000,
103'h3ce10f0b6c9f858c5c00000000,
103'h2273ac4384a05e585e00000000,
103'h02d5cd8ac2816d63ca5cd8ac20,
103'h1e858b6724f519a74e00000000,
103'h3cb054a826cae7321100000000,
103'h067aa375855072993600000001,
103'h14e5509b4000c7415c00000000,
103'h26d16b24c77b6ab6e200000000,
103'h1cb29f559c60bb522200000000,
103'h395ebab883322676ea00000000,
103'h1b5b48b49ee4c5cc86f5b48b49,
103'h3e589df2174380850800000000,
103'h28d15de6729ec939a600000000,
103'h2eaad92cf0f7672bbc00000000,
103'h36b67aea58c8c5122e00000000,
103'h1ca6e27446739e3f1e00000000,
103'h18daca833c2a19297600000000,
103'h08ad7bcbd8d0fb9dbc3ec02b32,
103'h2677944030abc620f800000000,
103'h1e0a71c6b85941ecd000000000,
103'h1b10ed8c60d0d62d02c43b6318,
103'h1541827b7edb47f3ba00000000,
103'h2443130858ec35801a00000000,
103'h26f069b62c2db7fb9800000000,
103'h22f70250d370cb03f200000000,
103'h3cce7118786134ba1e00000000,
103'h168127d3da58370af000000000,
103'h0920140f5926a8236a035e1619,
103'h26ecb8466ea7cff74400000000,
103'h192a278176c7e4069c00000000,
103'h02c8cb769cb49c4d0a8cb769c0,
103'h06bfa676b4dec3ce8000000001,
103'h24dd299a36a78f451e00000000,
103'h2ea27cb4fe6735bbd200000000,
103'h312fb3d663445f560a00000000,
103'h0e718744d0e6dc0b0830420000,
103'h20921e81c1168fe16a00000000,
103'h2a5a4503ce8817263a00000000,
103'h3289a141b11a35a7fd00000000,
103'h1cfd5cd59a747aabca00000000,
103'h1957f4748efe1bed7a00000000,
103'h14c91bf4eafb78c31600000000,
103'h1ec25a9b83536d37a400000000,
103'h1ad5ceea161c892c8e00d5ceea,
103'h315dbde476dee3c81200000000,
103'h14e3c8cc50b4b2b22800000000,
103'h23654c77401270969e00000000,
103'h353a3d59d4f63962ee00000000,
103'h1e2bb768f65b85da2e00000000,
103'h3cfc15402c95c3340200000000,
103'h2c8125c98ac17a9cfa00000000,
103'h1a18a6e986bd8fdd260000018a,
103'h1ea6616c733eb5a6b000000000,
103'h188fa1c98e575c903600000000,
103'h3f0ea55aacfdbdfcab00000000,
103'h2f4f2388c48d5fc63800000000,
103'h254d3194029c0520e400000000,
103'h0e89f545f0eb28a9a8449000d0,
103'h061e158815385a3daa00000001,
103'h2aaff3c6e4c24f839a00000000,
103'h12cf31cbeae0650bae00000000,
103'h3c8a74f1d69058d29300000000,
103'h1630e0c1695f8a9e7e00000000,
103'h070fa6cea6e9ff905400000000,
103'h18b0bc5f7c1ae051bc00000000,
103'h163236fc022a87206200000000,
103'h2b440a6b1cdb437fe000000000,
103'h28b56878b20d7a7be200000000,
103'h0b10c6169e5184e6fe00000001,
103'h2a8704064706ed5fb200000000,
103'h0e27c9165117b3765003c08b28,
103'h0ca3d1a63c9eb77c965ffbff5f,
103'h3f2d54b20ac68092e700000000,
103'h0e085ca4d66a52392204281001,
103'h24ea51f75697a6eb2c00000000,
103'h0ce3fac024a003900471fde812,
103'h2f7c5b058a8a55875a00000000,
103'h1cdb3bddd66e50477e00000000,
103'h20a46eef44eaab4d0800000000,
103'h3a0548ebe0c5e72ade00000000,
103'h38062678816a561a2400000000,
103'h0291598c7a6f9f060422b318f4,
103'h208adce7f575c57e8600000000,
103'h056f0b9076071f0b0000000001,
103'h0a192163d691fbf2f400000003,
103'h112d8d515c0107836a9642e6f9,
103'h10b19844e71a28e742cbb7aed2,
103'h06ab68b6f747b6389e00000001,
103'h30ac583406f94e7d8400000000,
103'h323f43a40ca4b7347b00000000,
103'h10d336977e510f68804113977f,
103'h148152723090530c8e00000000,
103'h0f772485836389a40cb1804200,
103'h1066451656e4dc163cc0b4800d,
103'h1efa1cdba65c009bbe00000000,
103'h2adf040976c245b21600000000,
103'h27543e43d4bc628dbc00000000,
103'h272d02223e9b66973200000000,
103'h3ceaa216e4efa4db0700000000,
103'h380442a74b1ca6fd4400000000,
103'h2ae028e9c60749142800000000,
103'h307871b9ff0b8bbb7400000000,
103'h34ac212168ebb4a53a00000000,
103'h1ccf7563d964265f3a00000000,
103'h100f70a38c104780a2ff949175,
103'h0d56b4f76adfbce47cefde7bbf,
103'h06a98506baef2d880800000001,
103'h28e809bb4645e27f7200000000,
103'h248ab4cf0cef67862e00000000,
103'h2f3da76376d771417400000000,
103'h20d056dc5b6226108200000000,
103'h0e5233dd489fcd73f80900a8a4,
103'h0519f35daa7024505200000001,
103'h06d11a6438c2582d9c00000000,
103'h3e5fb2ac3cdc4b8b4600000000,
103'h10507104c2ad65ef7ed1858aa2,
103'h2ce0fcd1410d189bbc00000000,
103'h32e1acee125d89a07f00000000,
103'h32a4b5387f3e8671c100000000,
103'h2f44090e3320335fd200000000,
103'h2c90c2d364c4e8985000000000,
103'h2cea95345208f1a68200000000,
103'h3ea1f135be99b479e700000000,
103'h1097d3a8ec8449ae3809c4fd5a,
103'h12ade97beb263ae3f800000000,
103'h3a88e7e73abe0e8ce400000000,
103'h336cd7f90e6bf808cf00000000,
103'h2aea7c84c8f4dff00a00000000,
103'h0eec6abebb61b7e9183011540c,
103'h1f1493dca74c346de000000000,
103'h28facb8774389f2c9a00000000,
103'h004cfb3b124d3309404d172229,
103'h20940adebb47fe90b600000000,
103'h3a3cd26b7a94f9cbc800000000,
103'h3c31ce661b2904aa8500000000,
103'h335f698d5665d715ff00000000,
103'h3ada37bdd297a57c1b00000000,
103'h3e9d047f04f70f097000000000,
103'h3ef4cb0bfed146c74300000000,
103'h197596437f6e4b464600000000,
103'h095c3890fc631652449f97615c,
103'h0ada805a94d8ac95c236a016a5,
103'h114fd72d9c34e526be8d79036f,
103'h149674c7e60f65815200000000,
103'h194b5da8765f3caeee00000000,
103'h16635cdb4af5b176d400000000,
103'h2a5408a3e2410f1f4a00000000,
103'h197999933aa46bfa9600000000,
103'h2eae9003e4f8749e7800000000,
103'h3842c3237c720e31b300000000,
103'h0ecca7b9ea209e3596004318c1,
103'h08979b6fa563615914fa7d1b58,
103'h3a06fb1ff2300912fe00000000,
103'h126ecf6ebac7a482a200000000,
103'h2748b1ef36ce9fa29600000000,
103'h254332a5483d6f115000000000,
103'h08a114b46e86210086139ada74,
103'h1e2effd692c953a5ce00000000,
103'h2e848f7b5a6a685a3c00000000,
103'h36a8bec2b8996830d000000000,
103'h050a5d1b681df7ac2a00000001,
103'h02f21c749ec6b66ee4e93c0000,
103'h12a32f73a2d1138a4c00000000,
103'h3cbeaacce4c32ffeeb00000000,
103'h20738e56f6665f728c00000000,
103'h2d46698d35250a3f7200000000,
103'h16dffb32549898966800000000,
103'h254aa061c2df02239c00000000,
103'h1678759018befd55f200000000,
103'h3e0caa30fd099db7b400000000,
103'h1cc5e91152821347cc00000000,
103'h0f17c088128ebd78ca03400401,
103'h03489a226e54a68a1c444dc000,
103'h0f387112bc6c67122e14308916,
103'h1931e5babeb501349c00000000,
103'h36ad6daa8ced72475800000000,
103'h24b7b313261f58021600000000,
103'h03169f05dcccc5aca40bb80000,
103'h1ae1f20ac08478bfca0387c82b,
103'h32624644429b17c5a700000000,
103'h16d00cc51e7d09d06600000000,
103'h215d2b4810df5014aa00000000,
103'h06b70f77a6af5cd9c800000000,
103'h2c956c67070c8821d800000000,
103'h170ee11c0cc397997e00000000,
103'h1e055fa1795904008400000000,
103'h36db2e3b9167e51c9000000000,
103'h346059af6e6d44be0800000000,
103'h38f20d45264872f99800000000,
103'h084758745aa8cca90877ca6ea9,
103'h12f5a7a4149ad9ee2e00000000,
103'h2a0bdbf05ce232628800000000,
103'h328f54faaed7da069d00000000,
103'h215b40fe9ae3b5f6fa00000000,
103'h2acff9ab8c730af1a800000000,
103'h06df8c46aece4bf04200000000,
103'h00d15144589e459bd0b7cb7014,
103'h2a9af0489f7dd1e27e00000000,
103'h2d484543e14f2326d600000000,
103'h3d68a530caea136f7400000000,
103'h3a57510df63258b35500000000,
103'h10e44286f49afde41e24a2516b,
103'h06ef05e26ef24ef21600000001,
103'h1b48ec64c0d691790afd23b193,
103'h3a8ce65686c5975b7800000000,
103'h100338fba00e83c038fa5a9db4,
103'h1a148984da9b6a16be00000000,
103'h121829002a9ea3126000000000,
103'h0cf259f484b32c973a79befbdf,
103'h0a92224458cb55976600000922,
103'h2b406e5464bdaf8bea00000000,
103'h268a247b2e4fd1d04200000000,
103'h0d727db45a904024a6f93eda7f,
103'h370e0384c11a649fd600000000,
103'h3b74deec8c8ce2543000000000,
103'h209969e0429ae5d8f000000000,
103'h360dc6a43d0fc4c57c00000000,
103'h2712638cdea92ea5be00000000,
103'h1631651554b6f549fc00000000,
103'h12dd48f1fcc958d6da00000000,
103'h122412a792fabdec2e00000000,
103'h0f7aa122a6d806de2a2c000111,
103'h297a5e4378fc1985be00000000,
103'h173110ae4776baa86400000000,
103'h02b11befeef118ebdc7dfdc000,
103'h002be51dc522299a22a7075bf3,
103'h247eb529c6d3458a1000000000,
103'h00cd9ebb86ff2aa7d4e664b1ad,
103'h229342f5ab7ddfd19c00000000,
103'h324a001baa4b7e8d2300000000,
103'h0622e6dbccdec182ce00000001,
103'h22cf1325fe28c19e7800000000,
103'h077a6a18074ba87a4600000000,
103'h14a3a0dba81abba04400000000,
103'h0c18562c6e9525b84a4ebbde37,
103'h126bcd000338c693f400000000,
103'h18e8057210511cc06200000000,
103'h22afe65e62bce9c06600000000,
103'h169282eafaa4ef327600000000,
103'h3b0a452fde54d590d800000000,
103'h20bace08b4e7587bd400000000,
103'h16bc73a1eef19dabb200000000,
103'h2e7b02fb8eac6bb46600000000,
103'h02de8187a568df5656061e9000,
103'h3496d5a494e3e251e400000000,
103'h1c36823d56c263d98a00000000,
103'h32c7cc81cd59397e1f00000000,
103'h1705827aa88fbbbb7400000000,
103'h20ac17c9da57883d4000000000,
103'h3e368f6af05d0ab7e800000000,
103'h34836ae592092281c200000000,
103'h34297fde513fb1ecb400000000,
103'h1e5f509284c31cd24600000000,
103'h20eca983faec9cb09600000000,
103'h14d70d2d594bed431c00000000,
103'h1aca9358793896c716000ca935,
103'h32fdcb704f0fa3f46f00000000,
103'h0ef4205a68da374ce668102430,
103'h24d711f51ad802bd3400000000,
103'h1205f0d2e8cc23179e00000000,
103'h386d6677cca3350cb900000000,
103'h2ee480111ea925dfa200000000,
103'h0d35d0f758168c576e9bee7bbf,
103'h055f249ac6fb0c688e00000001,
103'h27549b55d330dd5fe600000000,
103'h16ed471d969001faac00000000,
103'h252f18c4fee49d507e00000000,
103'h0a8776c3d4d1e46e140010eed8,
103'h36dae12b3800fd331200000000,
103'h355f28f2828873f6e600000000,
103'h097372b4786355221e8813cb33,
103'h1d6c59c6ecc27e14a000000000,
103'h023725477435f0c9182a3ba000,
103'h2202edfb10a24a900400000000,
103'h03572aa594d96fd77a40000000,
103'h1d0ebc7236dc5dd28a00000000,
103'h2088cc53783388781e00000000,
103'h1a38ccfdd44244ea540007199f,
103'h268b183836cb113dce00000000,
103'h04b6d34a1003de3ba200000000,
103'h1abeec2e768ef673d80005f761,
103'h28fa8d8afd45c9bdea00000000,
103'h0b7873d1d604b5ec600000bc39,
103'h24c16b567eff43775c00000000,
103'h0e0e4116c877b7493203008000,
103'h2eea0d4aec39229fb000000000,
103'h0c0ba33cfb4763b67aa7f1df7d,
103'h3f31ef1b6a3171016700000000,
103'h31577e71373d143e6200000000,
103'h2af4c510356f0359cc00000000,
103'h10cb2e4ee4c681cb02025641f1,
103'h32e8fb440ebb46db3700000000,
103'h3f38393aa086752a1d00000000,
103'h00c48b6f926f706e2a99fdeede,
103'h38bfe0fe52a7a9a8ca00000000,
103'h1481b858136c35185e00000000,
103'h3efed68d0b2c1616b000000000,
103'h0a0269ec1eadce6ec2009a7b07,
103'h29756db95eaca4fbce00000000,
103'h18901b2f68af0ee7ec00000000,
103'h1b16fdbdd0247ca14afc5bf6f7,
103'h28c9f662e8b497d0b200000000,
103'h162abd76c2cb958e8200000000,
103'h213829866c958bf16a00000000,
103'h14f4a47e02c049682e00000000,
103'h16d59c16e2f872ee9a00000000,
103'h026b2b8076ed176c9c700ec000,
103'h30cc50788ec2b3837e00000000,
103'h0ac30162112ddf03f60000000c,
103'h2779fbb3c0fa2f7c8400000000,
103'h252968f40abd30de9400000000,
103'h1ac5eda0f1372c92540018bdb4,
103'h1e2525d1556095865e00000000,
103'h32b23d05b12683274f00000000,
103'h063983b68e4ba8f8a200000001,
103'h257dfb4602fde5fe5200000000,
103'h32f99f67c93769b4e300000000,
103'h16d5d90feeb564fae400000000,
103'h28d895df60af0462ac00000000,
103'h0a26fba77684dd729a00009bee,
103'h2f73476de15d7351fc00000000,
103'h1cf6fce92a846ef97200000000,
103'h3730175f5af7b6675200000000,
103'h3318363836eeb3507f00000000,
103'h26853283ad1ecaafd800000000,
103'h394fa221213700e80e00000000,
103'h369e80b806bc336bba00000000,
103'h0ee515b63e0bd58cda008ac20d,
103'h1d1a5e04f6aa5644e000000000,
103'h186e7103848f6bfb2000000000,
103'h32f984ea22a9ca001700000000,
103'h1540cc3c7a183b039a00000000,
103'h3493e91bac11bfedbc00000000,
103'h0a915c3fc0528c2a3600000009,
103'h241e3b5ef4e67545e400000000,
103'h2254e47e3e77d185a400000000,
103'h18a3c8a124960ce49a00000000,
103'h3d046cb1c6eaf162d800000000,
103'h22b79cec9e8eba03fc00000000,
103'h3d51426d5c9326b5c200000000,
103'h1562b973bf4ac3a26200000000,
103'h130a3d5eba9c060fbe00000000,
103'h149cb2ac8efebf837c00000000,
103'h36bde1fe6108fce23600000000,
103'h35723805f6a5af8ec400000000,
103'h307151afed63918d2600000000,
103'h270c7169a2d5c9931c00000000,
103'h2ca650a6d2471b430800000000,
103'h13492cc63a538cacaa00000000,
103'h2e91b87466f9dd537e00000000,
103'h373dd5afb9430a19b800000000,
103'h22bfbc7e26d4c28e1e00000000,
103'h2088be8f9d12983dd600000000,
103'h18a54d4dbed254bbfc00000000,
103'h36bbb95f5e5b134b9800000000,
103'h0c152f8ab7006099588ab7cdff,
103'h084368442cbc19f8b67fb8de4d,
103'h2084393b78d149836e00000000,
103'h38975eeec014b1c79a00000000,
103'h310597eda298eb031400000000,
103'h1e743185da3049f1d400000000,
103'h389ee516ca35e1df7600000000,
103'h0c9ae22b28aa1365525d79b7bd,
103'h22ab91072248f87c1c00000000,
103'h18552ae62ee3daa74600000000,
103'h2a2f0eb7108f6bae6800000000,
103'h093ed4676ae4969496ed2179fe,
103'h0ef8ad7d1513a54ba80852a480,
103'h36fb7f0edd5279b31200000000,
103'h0ce22b47ea4b2730267597bbf7,
103'h3458432f6146a63f0400000000,
103'h06b2f1ab6e28d186ee00000000,
103'h2e214573228114b65000000000,
103'h32e212edeb340661bf00000000,
103'h20ee0798d8554bd4e000000000,
103'h3140a282ca375ec2ca00000000,
103'h2ebc0ef3aa25665ba200000000,
103'h10b8901adc6608de6c29439e38,
103'h1ae917a3cb2217d218000748bd,
103'h3e6eeb019adaa7ecf400000000,
103'h2b2c1d2236c3bf90be00000000,
103'h030eb59e7532aa925a59e74000,
103'h365756f91f5ec7b49000000000,
103'h36c21025e36d7d530400000000,
103'h1007713f98c4d44c22a14e79bb,
103'h201091ea0e86e4720400000000,
103'h244c5d26de8e55b19e00000000,
103'h06e6f0183e9ee79bac00000000,
103'h0cef005ca2eb44c28c77a26f57,
103'h2abbe4ed2ad234daca00000000,
103'h170fadefb6c135376e00000000,
103'h22f1cca3e17d1a249800000000,
103'h2e72d2f3b68cc8144e00000000,
103'h1cdf1e061b7e94b82e00000000,
103'h351d9df348f167abe400000000,
103'h031d5317e4d085b1fe00000000,
103'h309a226118ee23a54600000000,
103'h14a3b9be9a0b76bd2a00000000,
103'h152be5d44aa5991e4200000000,
103'h1aa57995de4952dcdc00014af3,
103'h06ef9309727538b12600000000,
103'h0927d0224f1ab247061eb132a4,
103'h276b83f8540a45507800000000,
103'h0c54d0ec9c321572c63b6aff6f,
103'h128770bdc29d996b1a00000000,
103'h0d2f494010f26a57b8ffb5abdc,
103'h12f1d4096279db157a00000000,
103'h2ebea4232ea924558a00000000,
103'h26bd89afc29af85eee00000000,
103'h215a08a770599c821c00000000,
103'h2ce8f1f6d6172631de00000000,
103'h1af1b65bb6712ed94e00f1b65b,
103'h36a39f16225a20d02400000000,
103'h16f0802f7d4bd72bdc00000000,
103'h2496fdcaf4ef7641fe00000000,
103'h0b54a1984adff6717c00000002,
103'h2683743eef76f43c7000000000,
103'h240c67b5b8cb95d4ba00000000,
103'h20e132585e4f0a13a800000000,
103'h10a5733d055b71c962a500b9d1,
103'h0a49aa93243ca421c024d54992,
103'h3564d625b6e2175ec400000000,
103'h164b978d012bc1f1ea00000000,
103'h16816307f4909817a000000000,
103'h1c12a04c4adc2fa4a000000000,
103'h06e081b2635d92ac9600000001,
103'h26907a773e7032f8e000000000,
103'h076c352e0450b4ab4200000000,
103'h1cd887fc6ae12f228000000000,
103'h3e210a6f704d64508400000000,
103'h00c71f8f0e25ec4cee7685edfe,
103'h02dd67a78d46f6bc60d3c60000,
103'h0644646b4d0e164b6e00000001,
103'h368c90518eeb7df2fa00000000,
103'h17222088562fe25e4600000000,
103'h04dd9d0c0cbc72afd600000000,
103'h3ee0104c22de93382d00000000,
103'h04f099d7a6bc30443800000000,
103'h1aeca156249c40905a0003b285,
103'h06188b32e88cda680000000001,
103'h3f00e7bf85797bbe2400000000,
103'h18c7d7844a9206f10c00000000,
103'h194af78d4a92eeb09000000000,
103'h3c6a5826a35ac634dd00000000,
103'h0b169327fca5bdc22600001169,
103'h1a3c49e7781015e8c801e24f3b,
103'h36f407980226a910c400000000,
103'h1d3eb3f91f62f2f83e00000000,
103'h26e4268f1456fa904000000000,
103'h2b2f56e73295ae895e00000000,
103'h288a9d281979d5187400000000,
103'h2a0c8c79c2a92bffa600000000,
103'h08f16ec3ad33c927bee153f209,
103'h3d2d4b9dd64055a18000000000,
103'h22fed7015e31c4652c00000000,
103'h214a377d5c5f10030200000000,
103'h223ec3f8ff5de7046200000000,
103'h0f67199c60a81e81be100c4010,
103'h12cfc4e142e6e27abc00000000,
103'h346a348b504dfc171c00000000,
103'h3263b438621dc0f85f00000000,
103'h2ebb1ae9d687f583b000000000,
103'h0cbaa01d08eba9bc127dd4de8d,
103'h2aa107caf8a6c4a5ea00000000,
103'h1ad56b90046164c2f200000035,
103'h2e27904d6e026c8dea00000000,
103'h1901aa8e8ad7d81dee00000000,
103'h0ac76e8bb8ff686b5e0000c76e,
103'h3733f72ed10112f9e800000000,
103'h2401e494dac88185a000000000,
103'h02d23e88d0fc78b47068000000,
103'h2b7a709ab6fe5d494a00000000,
103'h0a220b17f8d09bd21c00004416,
103'h3acab88f254b0c6cd300000000,
103'h063be78bee6d1784ca00000001,
103'h22a98f3d2a37d013ee00000000,
103'h35159437b173b79fde00000000,
103'h3f523504531d46dd0900000000,
103'h2ed9e23dc732db14b800000000,
103'h0ccea6fc048510190a67db7e87,
103'h14fb3bce335ef256d000000000,
103'h0c9b88403e2d9952d45fcca97f,
103'h16591b8f5328d5210800000000,
103'h264989f31ec45d614600000000,
103'h3abf086ff51d78f09b00000000,
103'h029379439a6702e3b8d0000000,
103'h0a95836a17260b53ae00000095,
103'h24c062b198b984974800000000,
103'h1caf9f5a624f08015e00000000,
103'h0abc54f3c70f6ab2f800000005,
103'h15300d70e4bf0a0d5a00000000,
103'h32c9d141af7b5f012300000000,
103'h2a1d19a9c2ab6c720600000000,
103'h06bf6a1336753db3b400000000,
103'h2871252fa092575d7800000000,
103'h2ee1ea596751c170ae00000000,
103'h22ce0e844ec2e6a04e00000000,
103'h1a659f213ca4d0f9b600000006,
103'h09726d71e072df7e04805907f2,
103'h1811931ffad87e9f4200000000,
103'h0f027a3ec54aec112281340800,
103'h12b647fddc5c7f311c00000000,
103'h150ee6b6aa5ef96fe000000000,
103'h36da64ed7c15416dbc00000000,
103'h157e61c3922428246600000000,
103'h346d4aaac8fe8d11e400000000,
103'h32b8b2c31d7ceed57700000000,
103'h1963144b52ea39803e00000000,
103'h3d22b74144a2ec435c00000000,
103'h3206825b9d06008eaf00000000,
103'h32e8da87db28b7cff300000000,
103'h0e4821898c2f3a2b8e041004c6,
103'h3c91a20b7e1814b36800000000,
103'h2e7e0ed0cd60363cf600000000,
103'h3c707c24c8f1d8487500000000,
103'h268ba148b76fe7194200000000,
103'h1cd6009834e0633e0a00000000,
103'h1138749b1b6c0486c2e6380a2c,
103'h12fb1edaf742051ef600000000,
103'h1eafa163477a79ba1000000000,
103'h20d40b04db7598950600000000,
103'h16d8d7e4782539f84c00000000,
103'h2749a94ad8f944fd2600000000,
103'h2cfc7fd02ed21ce19e00000000,
103'h3929d00f941bc62c7700000000,
103'h20ccb8e4001845fca400000000,
103'h3e94dbb0b842160c3900000000,
103'h3656437a980ecef03800000000,
103'h1ae9c82618a3aaa0f20000003a,
103'h149912fe0ef9ee1b8a00000000,
103'h0c60a3d2a8e3b641a271dbe9d5,
103'h3e6a4ab37c7cc93fb000000000,
103'h0a82c0848add6d125a00020b02,
103'h2c3ee0f68847b7c5d600000000,
103'h1ef4ef8412ca784a6000000000,
103'h388eb45341095940ea00000000,
103'h0ea542621efe48c4fc5220200e,
103'h30993d83568cfd183c00000000,
103'h1ad4f06a64323f7a5a000353c1,
103'h16db1b9bd4cb7cfdb000000000,
103'h14eaa00e2ea06d681600000000,
103'h2ef86d45867b8903ea00000000,
103'h209337951b6629121a00000000,
103'h3660415f095e9657a000000000,
103'h20f8c826a8f1cdecba00000000,
103'h3a31bc565e520f4bc200000000,
103'h1ae6398a014ad7726c000001cc,
103'h1400dfcfba7c93c8ca00000000,
103'h197a1c6d1662cd52ca00000000,
103'h04e526f72b63ad228600000000,
103'h0ea240cd02ddc98f9c40204680,
103'h1aaa321546c2f086c60aa32154,
103'h212eb72657653153ca00000000,
103'h3d16098a300f63691000000000,
103'h03610910903e1a8f6642400000,
103'h0c89d2268c542419966efb1fcf,
103'h1e758bc34eb52d2a2600000000,
103'h04c676b3dc3eff50b200000000,
103'h1d26c50d7ab48b140200000000,
103'h02c52df67f7b01c7de7d9f8000,
103'h36b7baf91aa1c6d55800000000,
103'h395f7525de66f4cbd700000000,
103'h17462ea3551eafc4f200000000,
103'h2ee17334cd7e24ead000000000,
103'h04f7b98e22c4538e2400000000,
103'h36afc6bcd0a5c6c2f000000000,
103'h06cec8b7549d80511200000000,
103'h2b0c7a76cd4d470de200000000,
103'h1ac85121121c0fc5360000000c,
103'h2d487b597e288a3c0200000000,
103'h0e6e6c54d8f0db5d1630242a08,
103'h0731dda1473956b69400000001,
103'h084295fb94a7c30b6c72ab787c,
103'h1e6f5e1b1ad9a0acb200000000,
103'h32c4b076a51c36a84900000000,
103'h200ade2f428b94c36200000000,
103'h128a629e7650453a0600000000,
103'h1ab1aa19175b23694a02c6a864,
103'h3eb2924068e58607c000000000,
103'h04cfb11004973020d600000000,
103'h0f7864a30249c2613e24201081,
103'h0e715d70061973714208a8b801,
103'h24c579a65691d8144400000000,
103'h24ff1be4650335844c00000000,
103'h26cfee434ac8af2aa200000000,
103'h2cea83036ec7cb0f0600000000,
103'h381e8b34d497b9525100000000,
103'h1ae46b7a80823c55be00000000,
103'h20ad814478a0c78a9400000000,
103'h323f4639128533051500000000,
103'h3098d63cb532b4498e00000000,
103'h048a1f92a671fa82a000000000,
103'h1afda53e560ad0bf54001fb4a7,
103'h2911f2749c94f051fa00000000,
103'h08ab72aff6929590521cf39fd2,
103'h1f77a734dea48804ee00000000,
103'h18b5d63c674ffab4e400000000,
103'h2afed60344c7a1e9c200000000,
103'h18dcc61c1e7d78262800000000,
103'h3c4d4bc5497c4e296f00000000,
103'h3f625973635914458d00000000,
103'h28c761d65ea6600ad400000000,
103'h16f40c231e08b97e3600000000,
103'h229e2e9606d01b549600000000,
103'h36c49f325cc42777b400000000,
103'h2f4424143f62560dba00000000,
103'h046a0900f526f5401600000000,
103'h3898a76be36b19545400000000,
103'h3297612b66d522554900000000,
103'h085a42629f6dc9c12c9bc5d1d9,
103'h1c7f79a790052aec9200000000,
103'h24cba62c995f6d4f3200000000,
103'h1082ec05f4dee6f6c2d2028799,
103'h250f54349aaa8d235c00000000,
103'h160986246a2d79295000000000,
103'h1808e300ce3ccd5dea00000000,
103'h3467ad2c654653825600000000,
103'h06a55e4ebe4f36832400000000,
103'h308d9c9472b6e3af8a00000000,
103'h06a35403795c41fe4800000001,
103'h2cf5d8d06ae9de92ba00000000,
103'h368eb11fb08d32963400000000,
103'h3e76bff21c830b669e00000000,
103'h3815b2741211bc864e00000000,
103'h2c10e6f450887c786c00000000,
103'h0af5fa074a9e2eec7e00000000,
103'h1a683fb076af15e0d000341fd8,
103'h075d90c042a50fe81a00000000,
103'h05649e565c0d4f989000000001,
103'h14f42864e26ae058d200000000,
103'h2e21e15fe6cf7eaf2e00000000,
103'h00feb03bbcc3a71410e12ba7e6,
103'h12808effaae58873f800000000,
103'h020fbd5c2ae438afb454000000,
103'h1309cc117e64c7af5e00000000,
103'h0ad359760174850b8a034d65d8,
103'h3e608dee937e511d0800000000,
103'h1ed34adb1f51aa930800000000,
103'h282a40775cb238819a00000000,
103'h30e5fdc2fa85835cb800000000,
103'h3816401a22afc3d41700000000,
103'h12c4d38e5295c1971000000000,
103'h0cc511958aac01b1347688dadf,
103'h2377881e5e70d53f8600000000,
103'h32af8203eb35e6d51300000000,
103'h26973fbd8cad6ef37000000000,
103'h2e14bf0e3f5cf0f75a00000000,
103'h013e401026f430b4e619386286,
103'h30d896519408efc32400000000,
103'h0aa8d36814472fd34a02a34da0,
103'h31267f72041fc624de00000000,
103'h15011c734ec8998cf200000000,
103'h20cfea297eef18fef600000000,
103'h3ea7a7a2d2f035724400000000,
103'h32c694ef72c01f9bc300000000,
103'h29054860f367c73e9600000000,
103'h2f0c955f642e5c2e0800000000,
103'h3002fb5ccc33a48efa00000000,
103'h06e996cc7a4039ee5e00000000,
103'h109051d7ed43354b2ca68e4660,
103'h0a9ed421f22ccc17a6000009ed,
103'h2adbb29a02bd1def9200000000,
103'h174c35a10f5bf2118600000000,
103'h3cfcf2967837a4ab8800000000,
103'h10f0e4d70e83da4c963685453c,
103'h1611a32f4a80cce30e00000000,
103'h1eef7f771a71b1ba1c00000000,
103'h36294dd0708354e96800000000,
103'h049ac0d55072d4608200000000,
103'h22900e26c69c2230f400000000,
103'h0a06285b4b36e3064400c50b69,
103'h0cedf449ecc6f12d0a77fab6f7,
103'h00591521f6cd19885493175525,
103'h05370a5a84bb0dd24200000001,
103'h0eb121c4041422f43808106200,
103'h25621c33ca4b2d4ebc00000000,
103'h26da07d098fc4f12c200000000,
103'h1e1f0cf5bd5e6b468c00000000,
103'h1c1f1fed223873172400000000,
103'h1f3355d8c357800ce200000000,
103'h2a92b9131e769ffa0400000000,
103'h0eee6b603ca9f5d2c65430a002,
103'h30a888f3e63caee5e400000000,
103'h369b199eb42b1a462000000000,
103'h3ce52a5666d3a33a0600000000,
103'h22a5db081d6ebcd8bc00000000,
103'h0210818c9953e72f228c980000,
103'h0ab7d6f6faf9c2373e00000000,
103'h068a46a77e0a43c3d600000000,
103'h2930599208c21abad200000000,
103'h274529554f4c61625000000000,
103'h3cade047b77cbaf45900000000,
103'h0f1059715cc1e449a600202082,
103'h1e7d165ed96fc4915c00000000,
103'h36abee0728801e02b800000000,
103'h1c272711c6fd34619000000000,
103'h391f1b10bea92268b900000000,
103'h30d8f3595ad0497a8000000000,
103'h0302903354ef648b3e00000000,
103'h3aac4b1004c857e49800000000,
103'h3a533a4e46cae817ec00000000,
103'h38a34bf543773327f200000000,
103'h12c3a716bcca6d763800000000,
103'h3ed366c3766db96b7b00000000,
103'h30ab7e54c93160823800000000,
103'h2a4e7dfe0704c745ae00000000,
103'h2568b0cf38b0459a7600000000,
103'h1d4d5116a2fec3987c00000000,
103'h0a9faac986677467b400000013,
103'h012364fea4b4c57e56ec153e7d,
103'h3eabe6796f547047de00000000,
103'h32e4ad8eb177d5468300000000,
103'h0b1c383c6e23bbbff00000008e,
103'h28bb3751e008694ea000000000,
103'h2a0efbe5aa24a18b0e00000000,
103'h1ab730c152dfd8dcf00000005b,
103'h3cd73ae37ceed4c29b00000000,
103'h0b1b00c598a60583ee0000011b,
103'h3b672ff6547d40676a00000000,
103'h16d800b21e98412d0200000000,
103'h0528aa4adaff71235600000001,
103'h2f6828a630d771d57600000000,
103'h334dac8575001c205100000000,
103'h08b070cc236844c680ec1a0551,
103'h3eab763fd4b5f14bf400000000,
103'h0ea5ecd6de666218161230080b,
103'h0e77d5435d11d857ec08e821a6,
103'h0349d9d02cb7c52eca9d9d02c0,
103'h1a8423237a2f9a722600000842,
103'h07745dc2be7974425200000000,
103'h10cafa7a18fd9765cee6b18a25,
103'h37336f895f71f5288c00000000,
103'h0b53a9c76f3cefa2a400002a75,
103'h18a37e77a5705f2c0200000000,
103'h246cc76a2ec408f37000000000,
103'h0833a7c28667876b142a1054c9,
103'h0a6c7d436ad44ed5440d8fa86d,
103'h3ae24266f207f697cb00000000,
103'h0ec866b67d7473db362031491a,
103'h127293f97656b6422800000000,
103'h1e8448a7871f1cf8a600000000,
103'h146a4c2ad891b0f21c00000000,
103'h3c584645f615f999a200000000,
103'h22bab43c4a8045c47c00000000,
103'h0173d874c8d88c0a7226323f9d,
103'h224c19a5ea934046be00000000,
103'h1eb60bc92b0718bb8600000000,
103'h1335f7860e5332617000000000,
103'h103629076d093e2a9c96756e68,
103'h160ee6933f3f35b0aa00000000,
103'h067ae465ce755eb81600000000,
103'h22edfaf3e484454b5600000000,
103'h0cb443e36cff29b1247fb5f9b6,
103'h2483cafd8eed24a50a00000000,
103'h3a9287c85ca168887600000000,
103'h1f16a34b402533860400000000,
103'h291f04197ab7bb4e6000000000,
103'h1e268e98d8ce5e99a000000000,
103'h251b3dbd42ed62b31a00000000,
103'h04b1556a2113f14bf400000000,
103'h266ca09d052f2f093600000000,
103'h00dfa71e4ae0847356e015c8d0,
103'h35210c39314d25105c00000000,
103'h2a4fd407312ccc2ea600000000,
103'h02928d21274dd867d634849800,
103'h1e047544509dac6f0600000000,
103'h0456e1dad23039902c00000000,
103'h1af67381b134aed47e00000000,
103'h20c2d157348b90af5000000000,
103'h0edd07948e8204310240020801,
103'h0c94ea40f044d588366a7fe47b,
103'h1d7d067d7f21dd1cc600000000,
103'h1e99d18e8ab6c75db600000000,
103'h16422d4ee733cddb3400000000,
103'h1d6c8d4046cd9f69be00000000,
103'h12dbc2b9dc0fccb8a400000000,
103'h076cd550387c59f8ea00000000,
103'h04b4af444a581cb2c600000000,
103'h2930571390c4f202fe00000000,
103'h15799e4c9479a1474800000000,
103'h1ad2b23e3ca9f85ad800069591,
103'h1aa82028d02396a76c00000150,
103'h22d5aac62cf648e5aa00000000,
103'h3cc82766869e690e7a00000000,
103'h2834454e287413d4a600000000,
103'h124a5b90a43c3b3b2c00000000,
103'h0e84087a8f7080895600000403,
103'h34b3fe4a20badc19fa00000000,
103'h22825d282e3ee4948800000000,
103'h38c4cfdae4f2e2deab00000000,
103'h33437dc8c6754006d900000000,
103'h3d32ac3ffe3a0fe1bc00000000,
103'h26dcb6d1307d8daa8200000000,
103'h3ec5a5f6ecb039ea8100000000,
103'h3ca177fb528cf0bbb200000000,
103'h3ef28a06925296b29f00000000,
103'h017dabf38ef40eadf238dd50c0,
103'h32865b8b0ce698b48500000000,
103'h103f450d0d6444a8126d80327d,
103'h02851f4abeeaa0331ed2af8000,
103'h071d903b1129e5402c00000001,
103'h18aa0fd952af048aea00000000,
103'h391d282c1acc94c5fb00000000,
103'h24f48526f376a49f4e00000000,
103'h0eb68254ea93cccb6849402034,
103'h0aa264c30e8851f25a00028993,
103'h193d4bbc1f3ed4474600000000,
103'h00a4c77b28e1390a54c30042be,
103'h1a82e7d9801e84c67200000020,
103'h20f4d50340c34c419a00000000,
103'h36ef141f5a46341b1a00000000,
103'h29282782bc3b091e5a00000000,
103'h054273f0732a1d3db600000000,
103'h1e7b45249b5244c07200000000,
103'h3a77629a5e94b8b0e400000000,
103'h30b9b42b3e0ffdd57e00000000,
103'h23370eda7887606fde00000000,
103'h06de86c76941149b1c00000001,
103'h04d84374cb7823759400000000,
103'h2366b8d31156aa3cfc00000000,
103'h3e052c06d52eedb1c600000000,
103'h132affaa7895a684d600000000,
103'h0e91e7e9369ad28baa48614491,
103'h1570f39d8ac5d2362200000000,
103'h2aa6a98ed957ba1f5a00000000,
103'h170b4d31eec8adbce400000000,
103'h38059759d86f574bbd00000000,
103'h129ab40d6e7aa47daa00000000,
103'h36f5a2f728803bd78400000000,
103'h34a84c003a1aefe4f200000000,
103'h1f23a2c6321092dc1a00000000,
103'h230e50d7e6b8dedc5600000000,
103'h1673a36744dc81a28800000000,
103'h315931ce28ead27a6e00000000,
103'h0759b019fe5e75e1b200000000,
103'h0e6ac141eeb7a7afda114080e5,
103'h3d34b146361157c9d800000000,
103'h30db22ed057c190bc800000000,
103'h0b6c670e42b0ca51fe00000001,
103'h255c2111328bed3f0200000000,
103'h2c0382c3fcf8544d4400000000,
103'h2abc3c40a054755e7600000000,
103'h2cf10ec90d57f8227400000000,
103'h32d6aba3761434631500000000,
103'h294835bce505432c2200000000,
103'h1cb2142396dbeecf9800000000,
103'h327067e8be24248c7d00000000,
103'h1486b3d05cd638b01200000000,
103'h2cb1341b0f46a098d200000000,
103'h2ae0f791e2cd54692e00000000,
103'h3ceca9d84f7e88843d00000000,
103'h0e1c80ab395f80161e0e40010c,
103'h3d22902e364c29ee6c00000000,
103'h386f404a0568aa99a600000000,
103'h168944cf028b3ac7dc00000000,
103'h0421d1d83afa7b11e000000001,
103'h2b19def79283bfe0e200000000,
103'h075e160556a591b91e00000000,
103'h270af7acc0bf70b0b000000000,
103'h0b43141c071d86b606143141c0,
103'h2875ab9d2d287e62c600000000,
103'h182c02ff376b927ecc00000000,
103'h1e87ec1a5ee13e1bf800000000,
103'h24a345e6370d411b3000000000,
103'h30dc266814952d358e00000000,
103'h283d854cb938731bc600000000,
103'h180a76b028149983da00000000,
103'h28b8a62f93521ed09400000000,
103'h2e7416ca2a5c9580bc00000000,
103'h08c4b49a52153bb04e68c7950e,
103'h1c4dc5864089527a7a00000000,
103'h1aeb6ff60a4e0714cc01d6dfec,
103'h28db3936669bcc9b0e00000000,
103'h222797f780873c911800000000,
103'h30893268ea6275c77e00000000,
103'h3e741f54cc8a0dbf0000000000,
103'h16ad13557d134027ea00000000,
103'h1481d3f13a875f7cb600000000,
103'h14ddd11e113472d23400000000,
103'h3e9c441266b646c36e00000000,
103'h36e4c4c5ba9417e18000000000,
103'h2b4085a0fb305bf3e600000000,
103'h1923a5f8f01520b9a000000000,
103'h193b39231a55a65a9a00000000,
103'h3e091310b2794c538a00000000,
103'h216b04dfccb48576a400000000,
103'h3afd52a2cabd98875900000000,
103'h06a4c11f6b289d672400000001,
103'h2aa1d5f6a625f009ee00000000,
103'h031837216ccab1295a7216c000,
103'h26431dc2d76c87200000000000,
103'h172b9ceb9a84be416c00000000,
103'h303cb97b80c7dc044200000000,
103'h3073c61556f378efdc00000000,
103'h1c7583d88730326b5e00000000,
103'h1ee3c8bbb6a3f880b400000000,
103'h3cd6cbe053197c593d00000000,
103'h1a91ab0932fd4514f200000024,
103'h0f400321eed410f546200010a3,
103'h0b1e8da60965bbfe7800000008,
103'h3ea110aad6a5bf206600000000,
103'h053d1008e2c44cc66e00000001,
103'h3cd6547be0655d714400000000,
103'h2343a9e424a26d7a2600000000,
103'h1116bb4ae078c1f6064efcaa6d,
103'h148f8bd202bc6bda2a00000000,
103'h3ccca91f92d327250b00000000,
103'h026f23de6662b2f70ce47bccc0,
103'h2eb40c17622f5c169e00000000,
103'h3971b646669e7ff50700000000,
103'h06ebcc4f94528c0c6800000000,
103'h2439097dccc44252ce00000000,
103'h2ae8f9a312b00ea26200000000,
103'h14c845def8e918203000000000,
103'h2246120fe2d211c34200000000,
103'h06166a4d369a57a23a00000001,
103'h36ab04dd5ae069b21e00000000,
103'h38efae0fe0f6d3ff5500000000,
103'h351d6f6296a1d8dcae00000000,
103'h121d42788e9186ec8e00000000,
103'h26b76d30c2aef64f2400000000,
103'h1632019b14cc38c7b400000000,
103'h24a36a04bc83a5f87600000000,
103'h0ab6ab4b12b5a7938c016d5696,
103'h3e5b737df75911984800000000,
103'h34af3200010fbce35a00000000,
103'h00cf2949be6b3061509d2cd587,
103'h0972c68bf51a62615234527553,
103'h22cc0b61b4e98bab1000000000,
103'h357e61cfbe5c52370400000000,
103'h0640752121285d98ba00000001,
103'h166db8d3d4a6bf687800000000,
103'h1cb55ee7dae734899800000000,
103'h16e690a6f354ed5d6e00000000,
103'h0f74149d0e0a4c454800020284,
103'h2729f62be4f0dcec3a00000000,
103'h148697233264f1894800000000,
103'h1eca6ca4188ee7b52c00000000,
103'h19632f826e157ed85e00000000,
103'h23063ea60cdfeb7c7800000000,
103'h0e9a2ab5e5431afee601055a72,
103'h2e93084f074959a4f200000000,
103'h271acd9d56e3845ad600000000,
103'h0cb811c405768ca9deff4ef6ef,
103'h3f3541672a915a473500000000,
103'h14f58c0937496c0b3800000000,
103'h32ff3050357ead726300000000,
103'h26ec58f20974397b9800000000,
103'h1f500e3dbd7369cbcc00000000,
103'h00451dd0a25fc2bdd45270473b,
103'h1883996ec2afd0fb9000000000,
103'h2440c27f42f4eecc3400000000,
103'h3b72250b5d78883af600000000,
103'h0a16f16340b94aba3800000000,
103'h3e1b8078fa2b6fc59400000000,
103'h34cfe08a47426128d600000000,
103'h2e792f67c45de1a1d000000000,
103'h029b06803a2dc22c161a00e800,
103'h19762852e8a6f193dc00000000,
103'h2a7cb9eb2b41f8141600000000,
103'h00c5acac44b82066febee689a1,
103'h1d6c810f2e34da522800000000,
103'h3241179e2efa86fe6d00000000,
103'h30bc9fc10c67080d9a00000000,
103'h1a7a1ff7fea81fabca01e87fdf,
103'h06efc095f164bf6cd600000001,
103'h229a3b860adedf64d400000000,
103'h2c3f3d7490ce9ffac400000000,
103'h024b4770b268db80ced1dc2c80,
103'h16ff71189ea818f56000000000,
103'h1c185a2d60f360661200000000,
103'h2b1022a6f8f2d17eb200000000,
103'h0ad68b1b540b2bac120035a2c6,
103'h1e05cf107e1b4e530a00000000,
103'h10dd2bfb0af1d96e5ef5a94656,
103'h22a7e94ba8f7a87ede00000000,
103'h2f65781af8d4d479e800000000,
103'h0c2e32965b7cbdc590bf5febed,
103'h2a123b64c8e235e08800000000,
103'h12e81da196106876e200000000,
103'h22b5a85d4122a3dbac00000000,
103'h2b580792d50ac17d4200000000,
103'h0e77248df6c069da8220104441,
103'h3b787769a218716d5600000000,
103'h3c8a32bc308f95fb4f00000000,
103'h3ebe91ea6b080d64f000000000,
103'h16fdb295e69240212000000000,
103'h24fd3d1be550d20b8a00000000,
103'h1415390f3b4e84a17000000000,
103'h34bccafdde4bc1bd5400000000,
103'h3e6c6a517360facc9000000000,
103'h2eae49c6261dc5ca6e00000000,
103'h0240fb46648a301be246640000,
103'h12223168123879e20800000000,
103'h034f2947177975286ec5800000,
103'h24dd1bf2a89ba6908000000000,
103'h2c88d468aaeacfd79600000000,
103'h1abebcfa8ec7ebca405f5e7d47,
103'h1d2d1f6e7c50c032ea00000000,
103'h3214f70ad70f7d2d7b00000000,
103'h32987537b33c9c9bf700000000,
103'h1f06c33c265193a6cc00000000,
103'h183cfd0ad8ea08de8000000000,
103'h0ec3f70c76f0cc1aa660620413,
103'h1a5a6e3b8e2dc9257e00000000,
103'h1a2d82069cf1c031f600000002,
103'h01522978784c2e6d84cf2bf2fe,
103'h0060d9c8d379b07422ed451e7a,
103'h37605633d4cbd9ec9a00000000,
103'h3a8d9bc4542cb3b56d00000000,
103'h1caca186ca8d09e94000000000,
103'h3617d5b6c41aa5ad9400000000,
103'h24fcba5ae2c747345e00000000,
103'h24ad78eb98df1ceb2400000000,
103'h3a8aeb31bcdbd7460600000000,
103'h18f56761228950319e00000000,
103'h3d7a893e1d143b635c00000000,
103'h02c6f24f7509a2c47e00000000,
103'h22f2784bf2842c029a00000000,
103'h3ef9d58e744b1e520f00000000,
103'h3c8a8302963d969e0000000000,
103'h162f6bda15376c2c7600000000,
103'h24ddf77610c1ef2f0c00000000,
103'h2610af14a6f15b092200000000,
103'h1c8e85054ccf527f3200000000,
103'h2949f193f2e00193da00000000,
103'h0b3cca4f0f6e869926000013cc,
103'h3ef1923936b8782d1900000000,
103'h1897b52c82f5427c2600000000,
103'h3f0d2a9f00e6d4b55d00000000,
103'h1762a1a5587e89e1de00000000,
103'h3d269f44d68bb480de00000000,
103'h18a315116cee56263600000000,
103'h3914cd5a2814f56b0d00000000,
103'h166d5a5840b80a7c7800000000,
103'h0e44713838ccd7d6a022288810,
103'h1aa73c99113a322ee2000029cf,
103'h14f85e201e7ea3671a00000000,
103'h345e75123825e0002a00000000,
103'h167c9680cc1e3e204800000000,
103'h33678fc6037cb3328300000000,
103'h1c8cbb3a18f949b34e00000000,
103'h26308a154a60d9795000000000,
103'h28fa38f0a8ed94b36a00000000,
103'h36e225ec4e1e1ec8b400000000,
103'h0946c61a761857b95caf48d195,
103'h32a4affbecfa7da5ab00000000,
103'h26637356b44143c02000000000,
103'h040fcb64e6e5f3bc0e00000001,
103'h2eda423bce496712c200000000,
103'h10bd10cc13593277aab1ef2a34,
103'h1e9a5d02013374b37800000000,
103'h20b8ecf810f0857f8a00000000,
103'h0abd70aa2e8ae2818a02f5c2a8,
103'h030b5b6f1143cf799c6de20000,
103'h0cb278ab9a014023ca59bc55ed,
103'h188d0a9b9e0c9b92da00000000,
103'h3458220b2abf143e7600000000,
103'h3eae1bfc434c1eda1400000000,
103'h1a47e566f6a440e53e00000000,
103'h10e2eef577525ce182c84909fa,
103'h248a9416d09a42487800000000,
103'h22f14d76a07d313dee00000000,
103'h24a425b08407c554be00000000,
103'h1efb3ecfa6f912cb5e00000000,
103'h0ca4b4d04c9d387be25ede7df7,
103'h0ce86d196a98774b8a7c3fadf5,
103'h2aa956a0773d2c1bd600000000,
103'h0e72057c432599354010009a20,
103'h1933c7236eceefd5b600000000,
103'h2e92c1467d40f551fa00000000,
103'h2e8a32b51574bc756800000000,
103'h24bed03f83077dbbe400000000,
103'h1f1906ff3091b070f800000000,
103'h06422d94955080b07a00000001,
103'h2aac497bf56987afaa00000000,
103'h228b21d8baabb5443e00000000,
103'h1d7177f16657fec03200000000,
103'h06e97e7b08e32098ee00000000,
103'h06b205b52754988a5400000001,
103'h38e4149eec3e17055c00000000,
103'h26c1d8ccf2f01cba8200000000,
103'h3af79bbb2cd431597100000000,
103'h18107f4252960a266200000000,
103'h1b7dfb53ce8da5e18eff7dfb53,
103'h0b298e6aa69e2523e200004a63,
103'h2ec53e3c011c2077b000000000,
103'h3d351f66cd45aee25700000000,
103'h1f3b0ab7fa0aed1e5600000000,
103'h0ece9beab6400c852220044011,
103'h25005241567b173d1c00000000,
103'h3c4e290fa549b327d500000000,
103'h1ee1aec04b4a05692a00000000,
103'h3c80218f46982e78cf00000000,
103'h105ea0e36479dd3918f261d526,
103'h3ab83774a0f9fec85e00000000,
103'h085b812db1589fabc4818f433a,
103'h2248d04fea10d7206400000000,
103'h00ce4deaf56c584e161d531c85,
103'h04cda8bf16b5289e0000000000,
103'h2ac7025b96837688f400000000,
103'h0118fba3dc511f480ab50d75f3,
103'h017bcc0c871821a3a249f6d814,
103'h374af4c347311d477e00000000,
103'h00cf461806ace95404be17b605,
103'h22d70df5bcf7de174a00000000,
103'h212ff51b7ec7242f5000000000,
103'h24a0fde4e09e32250e00000000,
103'h2f4323f5c2ce27408c00000000,
103'h0092335aa66f25256c80ac4009,
103'h0ed920d6d6b2491b2e48000903,
103'h1ae7328257447c75d6000e7328,
103'h06937652e51d9d4cac00000001,
103'h370de163ff04cfcf0200000000,
103'h0cf7719a84984621e67fbbddf3,
103'h38934aec3aa62785e500000000,
103'h3a73a0b3c69d99206800000000,
103'h207193c7ff30e40ca400000000,
103'h047456ab38a484c06a00000001,
103'h2c0f5fb0591618886a00000000,
103'h1050903b5c8a6f33a2e31083dd,
103'h3d2f59e6ca99cee3fc00000000,
103'h263f079edaea5f1f5800000000,
103'h08f33a175619b90622754188ba,
103'h04bd85183d58c0a4fe00000000,
103'h1f123f4cc64bfabc5400000000,
103'h0000c8654b097fd49285241cee,
103'h3ed9b09d291bbf215800000000,
103'h14cc51db2a1c8786a200000000,
103'h2617b3be28f63823cc00000000,
103'h3eaf105d7cc289fef600000000,
103'h204fecd162da3dbd1e00000000,
103'h2c0c8866a0894e1a9c00000000,
103'h22e5ab8282d93aebfe00000000,
103'h02b506c22ee5c352a061170000,
103'h1f46ec00d2cb6ed52200000000,
103'h1cb30efc948075975000000000,
103'h3ca88012f2c761982300000000,
103'h1e772c154e7a7094b600000000,
103'h312b9b6a4c22f0a7a800000000,
103'h12ab79946a9a1cbcf800000000,
103'h0aabcd55dac5b827441579aabb,
103'h337382af6e7131bbaf00000000,
103'h2ab5a89db91cff118a00000000,
103'h2e1abf33aa9081c0f800000000,
103'h1f19f28697462a5eb000000000,
103'h28dede00c460e9925a00000000,
103'h2014fb36a27adc18f000000000,
103'h1068177e0b59ba19b6872eb22a,
103'h2a4bb5866a6eb5505800000000,
103'h1c757ded7ad6ccce6400000000,
103'h13002fe6e6228254ce00000000,
103'h2b05bdf9429800424a00000000,
103'h0f650625549830293000001088,
103'h1e3303a1be9dee227200000000,
103'h28d7cdec8f02f447c600000000,
103'h189f1a8c2c35f7e98400000000,
103'h0afe676e140dc5d612003f99db,
103'h10f5e4792cace0623e24820b77,
103'h148b4fa6b6ab47d05200000000,
103'h2923af1c06a12c497e00000000,
103'h26f2067ada2c7bf03400000000,
103'h3ace23afc2502b0c3b00000000,
103'h39572146eb4231871600000000,
103'h2e8b66ae64105536d800000000,
103'h2860d85f5c67767dc200000000,
103'h3e62c6008af2dd2c2600000000,
103'h18b4deadf553b58b8400000000,
103'h1a4928e272b67b8c0e004928e2,
103'h02edc84dca6b5a3a02edc84dca,
103'h06f9de36e6b4831c7600000000,
103'h14f8d14c28a24b6a4000000000,
103'h194b79ecee9c29a12600000000,
103'h0e549e19c294faed4e0a4d04a1,
103'h0ec91c809ae074da3c600a400c,
103'h36f21e03e93512f40000000000,
103'h04bd6af178fe2f749a00000001,
103'h0324e1802ef04d788449c3005c,
103'h022152fc32adb869fc40000000,
103'h1cfe395274d299ea2a00000000,
103'h2010329cb6f3ece65c00000000,
103'h1d205b5b94f22638d200000000,
103'h0620d192f40258d58800000000,
103'h24cf00345222b4311c00000000,
103'h364fc8bfd94385c41200000000,
103'h3ec47e31bd1285f86400000000,
103'h1c2b59dc72624eb83c00000000,
103'h2e948e5cb326cce9fa00000000,
103'h1320770e0e5226c66c00000000,
103'h0eefe5837ce6b5231e7352818e,
103'h08d1d9f14e072c312c6b7ae031,
103'h36161d175cf711b4a800000000,
103'h14812d2766c8eba5f600000000,
103'h033e63fddcdf08bd54c7fbb800,
103'h2ae24ff7716035e4ba00000000,
103'h228d6822329e99e29600000000,
103'h372f92019e80e9da0600000000,
103'h309aa787010e51fc3a00000000,
103'h06e4c5c9b73de3fdd800000001,
103'h0c8f19f126d88b84d86fcdfaff,
103'h06d807fb2cbd514e8e00000000,
103'h1ea1dfdf394c6b3fb400000000,
103'h377a09bf8124733ae000000000,
103'h0490179d9ec6531a1800000001,
103'h397eb10096405cd99900000000,
103'h182a9bb21ad074773800000000,
103'h3322f1a3554f2577cf00000000,
103'h0a3fbacf6c79c129e8000001fd,
103'h0222d7159e9cb2cd3cc0000000,
103'h114650356adc6d9caa34f14c60,
103'h3a3a3dcc6cff44b24800000000,
103'h377d50db3e4594e7b200000000,
103'h213a2513f97fd2b42000000000,
103'h2a93ac19eefd238f5e00000000,
103'h1cc9a0bc913748a35600000000,
103'h3cfeda117acaf4bd4400000000,
103'h1a79a84e16949579d4000f3509,
103'h3174493ed4936f8b4e00000000,
103'h366c0dbeef0d17d96600000000,
103'h0a9b1ae2608161183a00000002,
103'h1a951cc316ed6ed728000004a8,
103'h0023b41da08889b988561eeb94,
103'h3a45bb037a1da67c9f00000000,
103'h2274d9c2bb415a9a4000000000,
103'h2c25599a3487159dba00000000,
103'h0ac34848d8fbef60760000000c,
103'h0ae9c0b1042148faaa000003a7,
103'h062ddf95cee491438200000001,
103'h3cb35914dace51f48700000000,
103'h26bfe831a0fc318a5600000000,
103'h2ac866aedcaf8a9f3000000000,
103'h30f22e26c36f72d0d000000000,
103'h060086e22d37d97fac00000001,
103'h36dd31921e2a07a66e00000000,
103'h06b60dcc652a8e889c00000001,
103'h333e74a5dd07c01abb00000000,
103'h22364e5022bdcde71e00000000,
103'h3f66017a16fc428cfb00000000,
103'h38bfbc4a793290dd1e00000000,
103'h174405a3769892573400000000,
103'h12d00f172f584ea1ac00000000,
103'h3019e672049c54452200000000,
103'h24600059d76c635c5000000000,
103'h10d8ab1ec68649ce542930a839,
103'h32e9e83aeae64a282d00000000,
103'h025373f8babef546f2ba000000,
103'h165953fbaca8dd81de00000000,
103'h02cb975aeefc517a98bad77000,
103'h36c424888755a5764600000000,
103'h14a2fbde48213cd13400000000,
103'h2c40c87afee56159ba00000000,
103'h3287729992885d380500000000,
103'h28ca6e32c0c925b30200000000,
103'h22630f423350984c9600000000,
103'h261ced22db1b067f5600000000,
103'h2abc2c5d3e7e15c18800000000,
103'h00e3c8cfa49b02e464bf65da04,
103'h16d48af50f572f41a200000000,
103'h1e15e5670e3af8114600000000,
103'h02724658650f83065619619000,
103'h254cbd0b4425686d6400000000,
103'h2cc236a28697aec5ca00000000,
103'h028edf7b6ce46bd10eb7dedb00,
103'h2696806598a6a2739400000000,
103'h30ada4561a3581ef0000000000,
103'h3eea30b400cc02549900000000,
103'h14be6bd7b279a6aab200000000,
103'h147712cc7163d75eb400000000,
103'h2ed65c34c52243366600000000,
103'h216b278c1a995602d600000000,
103'h14cbf538096fb2379c00000000,
103'h3aa6698ea8dad9c3b600000000,
103'h12e4b543fea6cefbbe00000000,
103'h2e45442fb84d388a6600000000,
103'h243f291e4a31edce6400000000,
103'h22a8c044797731fe1e00000000,
103'h08ed312e5cb65b1c682db5191a,
103'h2ed87113ff5f1b60e200000000,
103'h0d10e984084c4c8f3eae76c79f,
103'h357b4fc27724bda33e00000000,
103'h175ce7ff0335a7274600000000,
103'h16f4db57f6b0f6e9bc00000000,
103'h14ebea11cf0ddee8be00000000,
103'h1b2f455ae402ba40b4ffffffe5,
103'h16975e4738eea4528200000000,
103'h15351e5ad21de9ad6600000000,
103'h0883d55828b547f49e1b49565b,
103'h0ce06b3e3cea664f707537bfbe,
103'h323fbb65046e3ba79900000000,
103'h128dafde504ea6e5d400000000,
103'h02f98e05048e624adae0504000,
103'h1d1ab420561c12292a00000000,
103'h3026408b1815a02e2e00000000,
103'h0aa0089d7430544e84140113ae,
103'h37687795a75694d99e00000000,
103'h24bf48d8b0f69d771200000000,
103'h2a322c44e65f150cb800000000,
103'h08baafdf4d1e5de56ad2791d13,
103'h1b7387c836508a2a50ffb9c3e4,
103'h1482f48abe0b3a099c00000000,
103'h3e88fec4587ec1d1d300000000,
103'h0eee1e0aac01b65c90000b0440,
103'h2c719b366a8ab520ea00000000,
103'h3f45a28c7a78d32b9700000000,
103'h1124e3ec26ea6e62021d3ac512,
103'h3a82e71da53010ee7d00000000,
103'h10e2a0abb554f4daa2c6d5e889,
103'h12cd0f5aaed7dbf84600000000,
103'h0f30513540ba7ca3fc182810a0,
103'h307e0171d2878bfeaa00000000,
103'h38fbc29ce2b7dd33ea00000000,
103'h34ce78a29335dea5be00000000,
103'h1e790aa08b31a142a000000000,
103'h0ade19427e0019e53200000037,
103'h08cab3e31f792485bed9cbb350,
103'h296f2bb7a8573dc83c00000000,
103'h1b498231f021f1ab5afffd2608,
103'h195579eed8911d630200000000,
103'h16618b90f2da9f94f200000000,
103'h30e6c1b8cc301983ca00000000,
103'h34c335a8e291a514be00000000,
103'h26c19b44537866cd8a00000000,
103'h32511e42c73b9c766d00000000,
103'h30bb40d62efd37babe00000000,
103'h3b557ced614e55fd8700000000,
103'h26815e19510996d3b400000000,
103'h2525a612cb5f13c11400000000,
103'h2b058a82b0e071da6400000000,
103'h1ee2a6ad550617ed2e00000000,
103'h330e18d5810ba26fdf00000000,
103'h164321d15eee491d3200000000,
103'h04d73e8e52fc61f2b200000001,
103'h224bcd25a93f83c41200000000,
103'h16c673aa2f16c2526400000000,
103'h084cbc9e90628f780c1719f34e,
103'h1ac14eb0262903223a00000003,
103'h3f3242b47175bfc0cc00000000,
103'h0ce2ba7cca370e70f27bdf3e7d,
103'h06a9f4978a6951256200000000,
103'h12d3be2a574c0ba22e00000000,
103'h06268adf5cf60039b800000001,
103'h28ef175530c9be640e00000000,
103'h16eeb23bf6f049436a00000000,
103'h0e579e481edf60989a2b80040d,
103'h1d0c95f676ce12d49000000000,
103'h08b78dde8525b11cb0c91e611a,
103'h232c442aa33247132600000000,
103'h349143ba2ae9d4f1aa00000000,
103'h24d5a3e24c16191c4c00000000,
103'h0ae816df00a75cd6760000000e,
103'h34203af8657d00b8c400000000,
103'h028aa624ee651797c4154c49dc,
103'h38dee643248552902a00000000,
103'h3d493f7da60ff8b51800000000,
103'h025af58e9eeedef83cc0000000,
103'h2ce9ac585c381e75e200000000,
103'h04dd7ab9de9314048200000000,
103'h03569bab8b7cc05cdeeae28000,
103'h24dfb5524f5a3b16bc00000000,
103'h2657adf150b0d6c24600000000,
103'h0507c50636908c149400000001,
103'h004af01f9ce83a05e6999512c1,
103'h070adb95e2efff0c1c00000000,
103'h1c250222e23aef2bb800000000,
103'h02efff722a45cac19af722a000,
103'h1f4b88d6076acce47e00000000,
103'h168f4c3fc95acc56a800000000,
103'h32c30eb5a6a6552caf00000000,
103'h3031c0573d35a16c7600000000,
103'h18e63cba6ef8b0221c00000000,
103'h060586021e2a70795800000001,
103'h3c7f9ba07710ad33c900000000,
103'h18a0066b7c163335e600000000,
103'h30f612a2f895ced65e00000000,
103'h3844cefc9035d541da00000000,
103'h20bdfbcf832be7e4d400000000,
103'h3e47d5d63a70b6e16400000000,
103'h18e7e312da2eb2b0e600000000,
103'h2c1dbf25d97688872200000000,
103'h1289707ab25e6b99fc00000000,
103'h382109b45f7c2abfd600000000,
103'h1a2959cf71059b3a88014ace7b,
103'h19605c9b6a26a4eee600000000,
103'h2e0de7ee854ffebe5800000000,
103'h3619dedb9cb05b59c200000000,
103'h1ca200888abe43484600000000,
103'h342fbd7000d82223e400000000,
103'h36e41f465e7a22ac6e00000000,
103'h3ee87fdb12a9e01c7100000000,
103'h229d3bc98a8dff62ce00000000,
103'h11103b0048767f3de04cdde134,
103'h015b5c5aea13bb076ab78bb12a,
103'h0e20a061fa23f607b2105000d9,
103'h308fc4857c7f52629c00000000,
103'h1a8ce80bca9ff2c49800046740,
103'h0e008acffb2fb74a1400412508,
103'h2a87e89b96bc9f55de00000000,
103'h03333c6ee4bd2a25dac6ee4000,
103'h165de2a4cf4512c17000000000,
103'h37287b9f53784f305400000000,
103'h1022cbe3e8d631d522a64d0763,
103'h00d9bb7e5efead7474ec347969,
103'h144dd53eaf2179585e00000000,
103'h360701c06efb34d6bc00000000,
103'h2c387d7283490a156c00000000,
103'h0b402af9ba500bd5da000500ab,
103'h074685f5668889485e00000000,
103'h336e5a4970c8b4421900000000,
103'h0e916374370f3a377e00911a1b,
103'h2cfd76b46b7d9480ee00000000,
103'h04b995ca780ef7f52400000000,
103'h02fe3e28e40c6ea98e8f8a3900,
103'h310b9ac968c604740600000000,
103'h152831a16ac4429cea00000000,
103'h24c25cfa5acfdd665200000000,
103'h2a6b80486ef80f07bc00000000,
103'h1621124012ba6c021600000000,
103'h289ca8abbf25ec4a8600000000,
103'h26dc81b45446fe8a9800000000,
103'h3cec38233ce3a7365600000000,
103'h02f3fd99e2c028eaaa9e200000,
103'h1cb62f12a0ac610de800000000,
103'h329e4cd5e2a05ea7cb00000000,
103'h1ecd6923be568dba6a00000000,
103'h06e02ca7f2f4da904e00000001,
103'h10b31916d0c243b40cf86ab162,
103'h3d32669396a2705bfe00000000,
103'h0a5212b826558972ce005212b8,
103'h16c84c972287f0066400000000,
103'h163361066cda02be8c00000000,
103'h2560b929c4a24f55ae00000000,
103'h0b3081a91ad5b05c1c00026103,
103'h1655d39b3f366985e000000000,
103'h04031593c966eb2efa00000000,
103'h208a5a4adebcbeca3800000000,
103'h00b3ee57a4bfd45e02b9e15ad3,
103'h3ab332c0844a2ea8e100000000,
103'h34e8e0af46fe1d008400000000,
103'h368579cd00b14fc10a00000000,
103'h16ded1b4f49a30705000000000,
103'h1cf7fdfaea1faa3d5000000000,
103'h275b58e9c2fe7bf24600000000,
103'h36bcd0d91ef679ed3000000000,
103'h06cf98898451d2d6f200000000,
103'h0d7c90aa3a0ea3b010bf59dd1d,
103'h3e49330840de3c399400000000,
103'h311451588e5acce3ce00000000,
103'h02d5e9960ca3ffec10f4cb0600,
103'h16e954aa7cb851449e00000000,
103'h260b636efe8e3adaaa00000000,
103'h370bae6d16778f852600000000,
103'h1566c64efc82f2f42600000000,
103'h3f65de1cf28ea1613d00000000,
103'h251d472f86f567b03800000000,
103'h0b62eb1cc55b45cd2a0000058b,
103'h06201e8f29788cfcb000000001,
103'h3f6044f5b4db78197500000000,
103'h282f0cbd7afb96a89c00000000,
103'h18f33c357a5bdb9e5000000000,
103'h0c12b17aa28ae85bcc4d7cbdf7,
103'h2aaab3bc7d7e24914600000000,
103'h3a1e2e17c890d60be800000000,
103'h068d3f1bb23b89c86400000000,
103'h0d582bbdef59b7e02eacdffef7,
103'h36ae00bbf4e6f6fbe000000000,
103'h1a81fa4b423f22b9ce0081fa4b,
103'h08e6c9e678ed2375c405f549de,
103'h2a87234a136f1dc10600000000,
103'h3881348ddd55e7a77e00000000,
103'h3d623ccd86dd0af19000000000,
103'h028267c6fe5e3f7f6cdfc00000,
103'h008fb6363cc07c4cf2a8194197,
103'h120c22667f42e413f200000000,
103'h3ede763e40d29a4a2f00000000,
103'h328dd50792debcb0ad00000000,
103'h249b735050bd32eeec00000000,
103'h12698de6024b07f67e00000000,
103'h3e7a8c8fa6e67b46d000000000,
103'h2c5e25837850092cd200000000,
103'h2b207b27f8ca95bc7a00000000,
103'h3aa003bb6428bb3ff300000000,
103'h0e6a94454e493667ea240a22a5,
103'h091ba0160ae93a234ef94d1aa2,
103'h3b1cb5139953ce689e00000000,
103'h26e85fcda16f6e7ea800000000,
103'h34dcc5c79a8c23924000000000,
103'h121a62298174835fe000000000,
103'h3b4138aeb65149277a00000000,
103'h3abbdd9c896bab50fd00000000,
103'h1aa5f10904ace3ffb200000029,
103'h161c2807be68c19c3a00000000,
103'h1306e2665a0eb2a53e00000000,
103'h0542e5ec712adaacfe00000000,
103'h3eea94c38331bd135800000000,
103'h3f3f279a4774a2ffc800000000,
103'h3cfc7c0d455f37c34b00000000,
103'h14c88325829e5f5d9000000000,
103'h1cbf64eabe9adb6ad400000000,
103'h26e803c353635e905800000000,
103'h3685459bae22c37b1600000000,
103'h0a81bf37550ac73e6a00000206,
103'h221c98308a900cda1800000000,
103'h3b524c949711cc116f00000000,
103'h24eb5f88f82e6441f800000000,
103'h3ca735f87280b0d68e00000000,
103'h2a6dd3a6576c105f8800000000,
103'h24c47e2e54134657fa00000000,
103'h322cf4c7be8119fe5300000000,
103'h3ac3cfa32345982ca700000000,
103'h36db5b5516728cf46400000000,
103'h085ef76691365c9788b455f88c,
103'h2ef5d9d00711b7ec9e00000000,
103'h120dd637ce70af532e00000000,
103'h1a6b6acc3d6689233600000006,
103'h393b8c5510745f5b0500000000,
103'h28420a756adfca274200000000,
103'h1f5a4082651b567c5200000000,
103'h22e325e28c5d60f1bc00000000,
103'h24d29465eab7a1742000000000,
103'h363662444c9ac756ac00000000,
103'h3579fa49f26d5bbc9600000000,
103'h14d8e8cbe8a3be00e400000000,
103'h0295383f9d1db84ad6e0fe7000,
103'h1909292772f6a116be00000000,
103'h3d17e165f48bd9565c00000000,
103'h1293f5610c95027dce00000000,
103'h12b3c75d0aace3e3c200000000,
103'h2ef151a3dc40d944ce00000000,
103'h3c257d016ef4a0a1d900000000,
103'h3ee581b55ce5f245b600000000,
103'h0c3a88e7180b6f47241df7f39e,
103'h263c73fc96f0f0fc8200000000,
103'h1d7f3856e42b79e39a00000000,
103'h00b69d530b67ede0320f45999e,
103'h02d3f494e6e7263716d2539800,
103'h1efcbb1de69dc38a2000000000,
103'h111672a36b71b81f06d25d4232,
103'h275ba40c886e733cec00000000,
103'h0708c355d884e5e05600000000,
103'h0c9d08d63ee089ecde7ec4ff7f,
103'h38cf11e0c4e94d42b700000000,
103'h1172d30a50865618f4763e78ae,
103'h2e850770c85567f9b800000000,
103'h261c21b798c83b040800000000,
103'h1a93c5eb494d4274d20024f17a,
103'h14f4b761ae69642c6a00000000,
103'h1cdbfef108fd2a17b200000000,
103'h2e18ae7a1cf1e1796000000000,
103'h1b1d99073acde06a6afffffc76,
103'h0c6fc60928e68ee48677e776d7,
103'h2e2b5737820427ebc000000000,
103'h18e4127d9173edf4ea00000000,
103'h1e8eaf3cfe9f452c6c00000000,
103'h21072c66d68357a9fc00000000,
103'h0a663875341206e6fa00000001,
103'h36c96c6f5419334dd000000000,
103'h34a08e5e5f7f6bc30600000000,
103'h2f16f579d648d8325a00000000,
103'h0110b43f4ae96690bafd0d6802,
103'h061c79ebb9005c0a9000000001,
103'h204172e5f9111049da00000000,
103'h1ae5d7a33e2d8a3592003975e8,
103'h2ad31492e16efd1b8c00000000,
103'h04a9b8133a54d4beca00000000,
103'h1880b79e2627e951aa00000000,
103'h2468c772ead1a164e600000000,
103'h2e7e617d435259030c00000000,
103'h1a02f8a326bb2075f600000000,
103'h00dc6487d73981f33a0af33d88,
103'h0cddb9be303c7a96607efddf38,
103'h02b0b0597018df1e36c0000000,
103'h3cd5fff7bcf698dc6700000000,
103'h1eb6700bfea74935d600000000,
103'h14d062137c7d492d9200000000,
103'h3d26ceb15b33b9399300000000,
103'h12961a6d6f041b4d0e00000000,
103'h26fbff05eb2ae9fe6800000000,
103'h39092cd43ec1046bd700000000,
103'h0693a3d024bd0371c200000001,
103'h2f51d4059cc630460000000000,
103'h05141f882359d4162400000001,
103'h0701550910aba81bc000000000,
103'h06af8ef5d4bfc7a3e200000001,
103'h2b1acc545cc11cacf200000000,
103'h2a4c39f8e270aba2c600000000,
103'h0cd77bb38e8b77f7226fbffbd7,
103'h3e0e6589f8d7b1f00600000000,
103'h0705170446af2da39400000000,
103'h28bce52b84bd932d8c00000000,
103'h2ee55ef58ac2aa31d200000000,
103'h029950b6b57f8f5d5885b5a000,
103'h1024f467e264ee52e2e0030a80,
103'h235fc5bca6fe3f099600000000,
103'h3b582a3ef72333717b00000000,
103'h1e1338f31882f92e2000000000,
103'h354dd70494db236d1600000000,
103'h2eed6368f2ee5c602e00000000,
103'h0e8b2ed6e63c3364c204112261,
103'h254c2db6562996cdb400000000,
103'h149025c3e4b4c5a49c00000000,
103'h16af413e8b00f35af200000000,
103'h0cbcb9195e91191ed65edc8fef,
103'h28066458f4405a5d6000000000,
103'h1a79a66640fd1376be00000000,
103'h30a1ae18290377cfb400000000,
103'h12caa925027d1e35f400000000,
103'h1084bd50b51ecc4e1eb2f8814b,
103'h057f2bd9c6e975732000000001,
103'h3a76add9966e32c3d500000000,
103'h1971a7a91ced5e9d9a00000000,
103'h38e9bfae97640c773200000000,
103'h0e80a4022ed5b4204e40520007,
103'h2800fdc8e6bf73cee400000000,
103'h1aef8a53754017d112003be294,
103'h28cb757b9e411599f800000000,
103'h0c0b6d1af9309fed6e9dffffff,
103'h1f2118daa2fc15690c00000000,
103'h18f638692e0782840400000000,
103'h070b6fc8ce289b5ea600000000,
103'h1361bcc2671ed3c7d600000000,
103'h16e8a9a96d2a4390a400000000,
103'h3f6babf97e8c00530b00000000,
103'h14f630cd9574a9fc7600000000,
103'h38a9510052e055f5f500000000,
103'h027b44fae6d686c388da27d730,
103'h38777c861f7fd7c3dc00000000,
103'h2cffb46460fb1cbec200000000,
103'h34fc963f19729944e200000000,
103'h10d9ce0fc4724da94233c03341,
103'h148d8ca3fb6ee3e85c00000000,
103'h36c122fc0a48b1f82000000000,
103'h38efd612ded63e9c1a00000000,
103'h1491226e949761982600000000,
103'h36a4bc738e8737ab0400000000,
103'h10273a60e3185a199a877023a4,
103'h36f26a4658bd168d2800000000,
103'h3c93d8c7eae450ee0b00000000,
103'h16cca8e1a0d6bb346400000000,
103'h3e8cb0a65d6a93fc4e00000000,
103'h08651284b2373cddee29172cae,
103'h2cfa8af030c3ed844c00000000,
103'h3b745449ba290008fe00000000,
103'h2ac4d8d7a7238af93000000000,
103'h377ff161e297df42ea00000000,
103'h357246ca0c5cb81a9000000000,
103'h252889b682dca97c7200000000,
103'h0e07ccabf64ef0467e0360013b,
103'h210a9a9a9c7779fd0000000000,
103'h12a547cc2b7f46a8f800000000,
103'h129cad184a89e1439400000000,
103'h1370bbe0de2f290fbe00000000,
103'h0a93baeff0cbd6280a024eebbf,
103'h1e2e33fc033c9208e800000000,
103'h1f47f3b10ed04cf8d800000000,
103'h28eb94a9acfe80f4da00000000,
103'h10be5eb20a4674a5e83bf50611,
103'h285cfee27332094f9600000000,
103'h0238311bc2f06801a08de10000,
103'h2ce3b04deb4d66e41400000000,
103'h028db074ee8597ffd6c1d3b800,
103'h237e2541db69484dc200000000,
103'h36a0a35e5cf6f8c2b000000000,
103'h0eb3897c7f751e048a18840205,
103'h1113d67eb715c162e6ff0a8de8,
103'h00f9bb80c4c94adf64e1833014,
103'h0b48e8d094dd215e1a000523a3,
103'h308f0ee314d6dcdede00000000,
103'h154a52fa1e1fc5af7200000000,
103'h311b58740eaed4928600000000,
103'h0eb5a8cd62f9278ca458904610,
103'h022d1a84d2148000b2d2000000,
103'h097b691b22ca28ce16d8a0ea9a,
103'h2ee97d60e4f74352e800000000,
103'h200666392c72ac6e0a00000000,
103'h361c769e1a5c29ceee00000000,
103'h21470703bd6290081c00000000,
103'h2a3bc037727f06a63600000000,
103'h1a27bcbe12c60da9f200000009,
103'h368665b2bf01cde16600000000,
103'h2d41387658298a9f7800000000,
103'h215e9b420eaff0523600000000,
103'h06fb04b3faf128c88e00000000,
103'h3e5d7bcfda4fc40a9d00000000,
103'h36c1c0cd214ac8be9800000000,
103'h054f9069e0a8448e7200000001,
103'h228d5058d76a055b9400000000,
103'h3abc39105ab995c57500000000,
103'h2c3ae5d27d46e61e4a00000000,
103'h00045b5336031f2ea403bd40ed,
103'h35761562653e05012200000000,
103'h3e51d4cd244260545900000000,
103'h24e729fd5ab875b6bc00000000,
103'h06c3654bd90a4a83e200000001,
103'h1ea2bfc8fcf174813c00000000,
103'h1cc01f4742b4d9cd1400000000,
103'h3f1fdf19e35799961200000000,
103'h3b3814a33e17b8dd5400000000,
103'h0f5a94b07c3797f736094a581a,
103'h216e893ef66fac9a7400000000,
103'h3637579a84ca414af000000000,
103'h2d57bf8c2638ca89e600000000,
103'h228fe05b1d7022246c00000000,
103'h12ff992148c7e1b09200000000,
103'h3adefe81eb57c20baf00000000,
103'h2688a52d7e575b2cf600000000,
103'h396b1662f93659aee200000000,
103'h26bda9bcdebefedc6000000000,
103'h1cd81ec7572a153f5800000000,
103'h3f4a55dd7ce7befc3700000000,
103'h1e13e82098bfddc38c00000000,
103'h3713d412990a33a10800000000,
103'h2cd2bee0f61e1bc1a000000000,
103'h38bbbeeeae31efd43800000000,
103'h008c7df89b04aeb530c89656e5,
103'h231d1ac614c06da3de00000000,
103'h1ab7eb34944ceb9c7800000005,
103'h0a70d764b66a06628c00e1aec9,
103'h295bb3691321f1972200000000,
103'h224b3e229c92c8fbd800000000,
103'h2efb368006ee7c64ea00000000,
103'h10f81a79e939ba8788df2ff930,
103'h2a5f04d65734f1078e00000000,
103'h14e7e0c9e92d0b817600000000,
103'h1d0385b9528c1057cc00000000,
103'h2a0da70da673f121b400000000,
103'h215182e9847776db0600000000,
103'h2eca4fccee851de8ae00000000,
103'h23702831d0d6a0d23200000000,
103'h2aa210ee7ea0f09f2000000000,
103'h1847eacce01118d0f000000000,
103'h0a653b864ab329bf6e00000065,
103'h2a07aa2862fb148c5000000000,
103'h1c80b99cac6050129a00000000,
103'h0a9ab9b01967fa3afe00000000,
103'h1ac5d29474e8b3d7aa00000317,
103'h36a415383e836d87c200000000,
103'h357d6c685a49401c3600000000,
103'h1eb713ab10ed55547600000000,
103'h2358b528c56ac1bcd000000000,
103'h18e30a7e2321d567e000000000,
103'h0ef0cd5b457a8a90a438440802,
103'h1f47d0549e5d950ec600000000,
103'h3e8c28a26d4e626a0c00000000,
103'h233b42ad0c9632beaa00000000,
103'h2a0c321f8a225b611600000000,
103'h3757ac22ae5d9e0e2200000000,
103'h2100bb349969d02dae00000000,
103'h36f82cb08ec17c505c00000000,
103'h1a85d0eb2ec23784f400000010,
103'h0835d086e4ba64358247da59b3,
103'h24436e30bf403520b000000000,
103'h18badc08467605a79400000000,
103'h1af3c6302ab973d854001e78c6,
103'h0aeee7dd02744fe09a0003bb9f,
103'h1ea46dbf5d681610c600000000,
103'h329a28c26656fdedc900000000,
103'h0f05e96d06fb6bad2600b49683,
103'h142b1deff895946f8c00000000,
103'h1cc4a253869b7ddc9200000000,
103'h02c63cc7dac69bcc8cc798fb40,
103'h111ed529f88b3e201249cb84f3,
103'h2272d9393b517ae7ee00000000,
103'h2e5c71b80b705011e600000000,
103'h02e188136ee3294b2009b70000,
103'h302d3a3b5d3f9b032c00000000,
103'h16042a835f2123169a00000000,
103'h362c95b34e4e5d51f600000000,
103'h22c550f5255287d55600000000,
103'h3d4135821c7f1d88a400000000,
103'h34fcb5123f446e7dca00000000,
103'h0ad957b8fc85a3ffe600000d95,
103'h2f0457b1b08259122400000000,
103'h3881df7fba5bb0cb2000000000,
103'h1e7e84d66860087cd000000000,
103'h04bf98aae2e1e7fc8a00000001,
103'h2486507f41606cd2f400000000,
103'h36cf6165c520057dd600000000,
103'h017423176aa655fd160d3c8a40,
103'h3578ed45e175b762dc00000000,
103'h0a5f9f70e0e9da7a4605f9f70e,
103'h22a6be6ed762c7c02600000000,
103'h3e0de2eaa0c267310600000000,
103'h041b5d638269259fdc00000001,
103'h2a9e8f3f4177088a7e00000000,
103'h300b9b95449265ee0000000000,
103'h0edb6fab6f30f52d42083294a1,
103'h0d6daaf2a03c90c286bedd7953,
103'h0d690bd9af18006df6bc85feff,
103'h0edb754b3a85ab60964090a009,
103'h16e044aac6eeb73a4400000000,
103'h0d16093796ca2c857eef16dbff,
103'h22885e86ecaa71304400000000,
103'h2712b44438c07a67da00000000,
103'h2522b5621a48d8eec600000000,
103'h29216dba405b8d32fe00000000,
103'h04ea5297e47e42951800000000,
103'h0a5da8a5cc9fb04f580002ed45,
103'h0a91791b908a02e73c00000001,
103'h230e22801ce7ab8d0a00000000,
103'h3ce65917a67924a89a00000000,
103'h383cd24448874728b700000000,
103'h0232fbc0446da0405c78088000,
103'h1eb328237eaa7284a600000000,
103'h141b0013c0dd6e44ea00000000,
103'h32fbfcac9e9096686900000000,
103'h1964406e34ab967c2a00000000,
103'h033a247026a79328c8d1238130,
103'h2cba7af6be0bd396fc00000000,
103'h16183fc24045f8072200000000,
103'h1e069af62c0072fde000000000,
103'h1ca08ca64318b2c02200000000,
103'h3ee2117f221f4db64f00000000,
103'h212f69eefebfda5c9200000000,
103'h02c2ba65fca1ebdbb4f8000000,
103'h10567ddadcd155cab2c2940815,
103'h2202f40fde941030ae00000000,
103'h16ceb7fb30ea8e0b8c00000000,
103'h085a564312ed821b6a5bea2c3c,
103'h3887e066aabc3a169b00000000,
103'h0486c054f3169059ae00000000,
103'h2e19b073ea9e70c05800000000,
103'h0a972e9e6e2531154a025cba79,
103'h39022ee45f3ee1893700000000,
103'h11296940e8d61027a429ac8ca2,
103'h1b6733f720d83f0c02d9ccfdc8,
103'h11436f6db001a84ceaa0e39063,
103'h3644dbf98a68dc440a00000000,
103'h38852a0e9cac4bb1bb00000000,
103'h249b884b52f127ab4600000000,
103'h2e8a25940b7651b9e200000000,
103'h2a7a6b29af11da053400000000,
103'h30d38d035e9bff993e00000000,
103'h12d8fa8ec9166ac2ee00000000,
103'h06cf8fc578e9f7c64c00000001,
103'h053c76b60ac2f2551400000001,
103'h32bb37abd092821a8d00000000,
103'h3ed5f83ad4cef8d09700000000,
103'h1307238cc88a307c6600000000,
103'h1e2246a5066028b73a00000000,
103'h35005c125a674c440200000000,
103'h1a70f39a388992e90a01c3ce68,
103'h16b083f2ae89eefb6400000000,
103'h187a44c788fae2959c00000000,
103'h22a42e539eab66884a00000000,
103'h07356423b925ab4fd400000000,
103'h24502cdcdac9d9a37200000000,
103'h2ef4e49162ff3dc72a00000000,
103'h02947edb874f6aa40651fb6e18,
103'h36df7fadf5444f356800000000,
103'h21502bd038d8ce10ee00000000,
103'h268ab195eeb84dbee200000000,
103'h0ec47522ce08798f1a00388105,
103'h3d4da353b6932b250800000000,
103'h201b20ba0557a047d800000000,
103'h3ac16c3142a5439b8f00000000,
103'h0520056762c064559200000001,
103'h1c87182c9c81d086d400000000,
103'h2a815616e0a1d5ee3600000000,
103'h3cd33448fd28ee1ad500000000,
103'h12ca5616a6aa4431b400000000,
103'h0881dc39e57d787ab2fe5221ab,
103'h1cbb32e3f647ce915800000000,
103'h12965f7c3ec9aacb3c00000000,
103'h049a7a2f5c84ddaf3200000000,
103'h1d48d9142f1b3d2b7200000000,
103'h1b74b073b2b5b75aceff74b073,
103'h0ce856648efe906efc7f6b377f,
103'h3e25a720a97340e2ae00000000,
103'h0ce7d58bf65b97473c7febe7ff,
103'h08c54122b4813e67e6223fa2a9,
103'h37586414436913f3dc00000000,
103'h34ea1774ca2e55169000000000,
103'h1aef0bb80286b92ad2003bc2ee,
103'h374f97427770d09f9e00000000,
103'h07316134d15fdc57a000000001,
103'h1b7c3f1b06af739a16fff7c3f1,
103'h38f57217cce0d4cee600000000,
103'h18f55e3f675d13e9ec00000000,
103'h2e661b069e528601b800000000,
103'h1436b4257747e4412000000000,
103'h00b6c0de64adff47beb2601311,
103'h3817a26638e4b36d3700000000,
103'h18d597d7f89b744b9a00000000,
103'h18e6134b72b316b1d400000000,
103'h0e3e73000a88ae89cc04110004,
103'h2844d1fc626ec1d53e00000000,
103'h3c2fe465f0ad34d54b00000000,
103'h0ab66b1b1af206d1ac0000016c,
103'h08f008821721eb379ee8f1dac4,
103'h12b25472e0d85652b800000000,
103'h00e36238eac85ed4ced5e086dc,
103'h1ec1a4d43d7ab347b000000000,
103'h1691ee413d5e15809a00000000,
103'h248422e5da1fba54d600000000,
103'h144eaddd30b1a8961400000000,
103'h2ee197a95635cb7bee00000000,
103'h06ef34bd2a8479592000000000,
103'h1b5ae7519b66110276fffffff5,
103'h08e6543ae05545bfa05988c2a0,
103'h292369ba3ab02d113a00000000,
103'h1e964ab58296814c1a00000000,
103'h008da509ecb9eb0654a3c80820,
103'h3aeb1060cb5035bbd900000000,
103'h169dc1774adddac5c400000000,
103'h2b009f9f06c8eb268e00000000,
103'h02f9ff12dd66ac9ddaf12dc000,
103'h06ad498d07674c3ce000000001,
103'h16b0c9c30b614b4fbc00000000,
103'h309224bed00e94dcc200000000,
103'h103c6ae126bf5e9fccbe8620ad,
103'h0c4d5da15751835e9eaeefffef,
103'h0ec59c9e668dee3fc442c60f22,
103'h1c9f26eb32db4be11c00000000,
103'h3a874614c2a0e87f8200000000,
103'h3f2ec3de1f400f6ab600000000,
103'h1b27c50618c7557f78fffffff9,
103'h1eaeb46dd6f6195d9600000000,
103'h1510efb6b31dde63ae00000000,
103'h0d14137f10cc92d184ee49ffca,
103'h235746b224dd82883600000000,
103'h1161cf64b0f1960746381caeb5,
103'h15627174d248dcb96a00000000,
103'h0c80f1e8a2aaac1e1a557eff5d,
103'h126c052df60d1d92ec00000000,
103'h3e349afb828e0f7b8e00000000,
103'h18eec6d056fa14a98600000000,
103'h06f1cf5e942eafa50800000000,
103'h149f840aec1d76755e00000000,
103'h1a5a564a320f45d3f200000016,
103'h24a3380508aec9dee000000000,
103'h02e62e6962092029122e696200,
103'h3657d472c6ac582e1a00000000,
103'h16e6f0f18a9286977e00000000,
103'h2885534440ea5b0a4400000000,
103'h04d27f75d6d14bfbce00000000,
103'h0228cbd07e569f400e32f41f80,
103'h062b705942291eb5e400000000,
103'h16c09b798551ea866400000000,
103'h254021a40c7d5adfa600000000,
103'h0a90f3ca633df6592c00000121,
103'h2e386530c77e17fd3800000000,
103'h1408f54d110f0bc79a00000000,
103'h002b6fefbe4770f8603970740f,
103'h38cb4572155066457200000000,
103'h12a9114d947bd6353000000000,
103'h3504f5264e471ba74400000000,
103'h266fe4c6a0f02cf4da00000000,
103'h1622455f54f5221b2800000000,
103'h1c250c3d7a6506e1c800000000,
103'h36a3a950d2874c411e00000000,
103'h1f69620b6eac587e9800000000,
103'h271f47bae45001cf6a00000000,
103'h04ca4f8582b963dad800000000,
103'h1eda5e31e8d8ab95bc00000000,
103'h0971b91f6ea2fb1b3ee9a10228,
103'h22b56c8b8d7d594d2800000000,
103'h1e4921c714ef126c9600000000,
103'h1e963add76a47ef82200000000,
103'h06bbff8996eda0bf3600000001,
103'h1c84bf50f483db9cae00000000,
103'h3ecad8657b3fdb264400000000,
103'h350003e696c49a773800000000,
103'h22d9ae5fd48f72dcb200000000,
103'h26a0f998488f76c34800000000,
103'h1eec206d6d6925231c00000000,
103'h10772268d20a1ebb643681d6b7,
103'h18c6bedb72f63f28d000000000,
103'h34a5ce2ac36d6191a400000000,
103'h1b14543d5d34206d16fff14543,
103'h2aebff7310d9ee97d800000000,
103'h0ecdc9642aee42d53466202210,
103'h24a5d27e16da42484600000000,
103'h3eeb3d29a4a80bac7100000000,
103'h3364c8424a4dde2a8700000000,
103'h38b841f2c9391b542c00000000,
103'h2af9fe787a9de3967600000000,
103'h3115fd46755625893e00000000,
103'h1cda07c0de502401b800000000,
103'h12ebf065ce6621482c00000000,
103'h1136f45eec4029090a7b65aaf1,
103'h0a1fdbee7f2c196eda00007f6f,
103'h375ee90751630dcdc600000000,
103'h02ee1a21da82e9bc44dc3443b4,
103'h1ce36c8490e1d2c39400000000,
103'h2218e7f052cfece56e00000000,
103'h267a7ccaeeb3596a0000000000,
103'h3c3f1f7350cc415a5300000000,
103'h2a86abd7f946be254200000000,
103'h2ab00b003485dd989200000000,
103'h3ea9570dde0c89708b00000000,
103'h0155fc858abc9470be09487b24,
103'h12cee3578965eb7e9e00000000,
103'h1e8e884ec8bbe8042800000000,
103'h1cd40ade9a8acb5bb000000000,
103'h3a2616def91953aa7900000000,
103'h2334b75016ed5e891200000000,
103'h12a9433fd11375680c00000000,
103'h0ad9b733b5482cb8220000366d,
103'h1e94f68346f16ff7f200000000,
103'h2b69897d52cb272ba600000000,
103'h0d2b7b0071601daeeeb5bfd77f,
103'h3f00e1eb9ac9a72c4100000000,
103'h271e758ee6f5222cb000000000,
103'h142d792a24f604184a00000000,
103'h1407a3f10b1479a73000000000,
103'h0441ec66de41f2d15400000001,
103'h0e45dc08f34996c26020ca0030,
103'h3e3eedd7b68b83293e00000000,
103'h122e03bec4d15f323200000000,
103'h3231934d02104d09e900000000,
103'h337715ac973e50c8af00000000,
103'h24062ece886fe415b000000000,
103'h0c20cb19bae6f9c246737dedff,
103'h3a0cc6971eed2890d000000000,
103'h2d090f1e6c0df3aa8a00000000,
103'h3243a86e671aba41ab00000000,
103'h02ee25d41323c9601697504800,
103'h0f7f9cfc066771ce7c33886602,
103'h38fe3cb4c95597a29000000000,
103'h0e8ad01816d5349e9640080c0b,
103'h0a321dbd0ed371535e0000321d,
103'h1afd34c21d5e416b760000000f,
103'h312fbd95a8905f288400000000,
103'h10b7de0bc28d93eaa215251090,
103'h0715332074bd51804a00000000,
103'h0b45f98884752f8c0c028bf311,
103'h2cd5015c0a8a62ac8000000000,
103'h36f4685814d05c350400000000,
103'h04a1633ec2a55d910e00000001,
103'h040bafa5b899c5e92400000001,
103'h0aeb2b98bd3b2927e600000eb2,
103'h19550a384246d8cd9e00000000,
103'h3c8f450ccd3204665d00000000,
103'h226edd7264870e9e9e00000000,
103'h02e83bc1231653ab6a12200000,
103'h1e9cc337c485311dce00000000,
103'h3c98237c066d6cdef000000000,
103'h26c58826a50a3016b600000000,
103'h3479fb6fe0a25392bc00000000,
103'h2644c2648767dbb96200000000,
103'h1c94ba76fce1d7294200000000,
103'h19521f686326998dca00000000,
103'h3b19b4707ebb5404c600000000,
103'h3e839d0b570d736d2800000000,
103'h0955615f932727dda63923411a,
103'h0f08fcdd10aac4e8fc04626408,
103'h36e331e8580026488e00000000,
103'h1d78baf8660923259e00000000,
103'h191bb7759cec550df600000000,
103'h28e5dbd0786510065c00000000,
103'h065ac5145080c77bf800000001,
103'h3ecfd4a0b866a34c7100000000,
103'h1b4e0752c0c16860c2d381d4b0,
103'h14b88f12be913d017a00000000,
103'h048826d918df44543a00000001,
103'h06d8861b6c97d366f800000000,
103'h028f88aa331ffa401288aa3200,
103'h3c07f399b8f8805b7f00000000,
103'h36119b8aba880905b000000000,
103'h08fa87cff88ffc9f6a3abda849,
103'h077b477c2ea1982a2400000000,
103'h391c0168769c1ffa1d00000000,
103'h22b53bb03c1767764a00000000,
103'h06d67efdb43368dec000000000,
103'h2487beea96e8a48efe00000000,
103'h2eda97019ebf238cb200000000,
103'h30c98f12c346e2774a00000000,
103'h2ecfee9a31217978e800000000,
103'h2009b70060eb088baa00000000,
103'h2a2c23f58ebaf725da00000000,
103'h130db47770c4ae263c00000000,
103'h3c3627709af0d21bcb00000000,
103'h188013e2aefe86933a00000000,
103'h14b508e06b34ae03d600000000,
103'h1ea4f50402b4c1e68400000000,
103'h1a598f4dd669cac6ee00000059,
103'h30fefbb3770ebfcaf200000000,
103'h34a2eeac50684f18c800000000,
103'h237b8fa900674acc3e00000000,
103'h1508f28c340a39788e00000000,
103'h1e0020365685c9218e00000000,
103'h1d060dab6c8ebbadc200000000,
103'h2d744a394a8edbe41a00000000,
103'h3a49d1936694e98f8600000000,
103'h3e299266130933c8d000000000,
103'h188f1c5a4e53055c3600000000,
103'h1e8361fc4d7c97c24a00000000,
103'h2f068382650bb41c9800000000,
103'h251e8e98028f1618e400000000,
103'h2f3fcd767095999b4800000000,
103'h06b411b114b428334a00000001,
103'h2aa4edae04f3f5a9ba00000000,
103'h32a17dc78aa8075acf00000000,
103'h3d2d23f9f64cf508d200000000,
103'h364e63c7a8ee72d05e00000000,
103'h0723cbc8a71b96ca5400000000,
103'h18ed29735c69fa91fc00000000,
103'h365e8e78e28dc65aa200000000,
103'h0b1ce8873d7aefce008e74439e,
103'h08c9b565f2d97e46e208659188,
103'h2a92190efef666ce1e00000000,
103'h2ac4774a06c01c341200000000,
103'h0e849bdfb1523543100008a188,
103'h2cbfb0435d16ac8d1600000000,
103'h3ed442edea9b486cc700000000,
103'h0edf3c66965af8b0222d1c1001,
103'h24aa5213562f3b9e0c00000000,
103'h2cc79d03250e7804a400000000,
103'h0efb94800ab8ca17fa5c400005,
103'h1ccad469b680671b1e00000000,
103'h00f50d03847bfb9b28b8844f56,
103'h3a4e813b6046d004df00000000,
103'h18b66d77e13bdd086400000000,
103'h02d723cc5a8a5e43c4ae4798b4,
103'h2178413bf540cbbba600000000,
103'h04955a46b617ef880000000000,
103'h0af94356569030c3f40000001f,
103'h3099096e5c258b0aaa00000000,
103'h30c32dca271ece610200000000,
103'h272e1de196b7d7cf5e00000000,
103'h10b0fd81077b0599849afbf3c1,
103'h12c40de46ca9237b1a00000000,
103'h30fca9527e5a20fc2000000000,
103'h34541321911e2ee08e00000000,
103'h0f6354c0031ad8330c81280000,
103'h30ed9bf7f66eeb549c00000000,
103'h3f2106ab06d240149f00000000,
103'h0aae925a36bfdc0c96000ae925,
103'h275a4ce9f4e0e2b79c00000000,
103'h0720dfacbe8f7511d200000000,
103'h1c565dc424e9c1fbc600000000,
103'h385e1bf02b0aa1a88400000000,
103'h0a25b628c660ff6ca80000012d,
103'h10ce3318febf1b5cd4078bde15,
103'h1406251b08e4d1859a00000000,
103'h3c27d918d8b3049e9b00000000,
103'h10542ebf2cb929b9a2cd8282c5,
103'h2ce183d22ae102d27c00000000,
103'h062df441fa353191a800000001,
103'h285f36376616b563d200000000,
103'h24437ccb6d44a9a5ce00000000,
103'h0ee0ed1916a3dfdd3450668c8a,
103'h205f60393ae75ca8a200000000,
103'h2e1304eb08c849c1b800000000,
103'h24dd5f00aa27a9faf200000000,
103'h06ec62bc193aaee5fc00000001,
103'h3e9f4654bd180de6a600000000,
103'h30398696020470a2be00000000,
103'h2c9c109900a3b6f77c00000000,
103'h13264496f2dd3d8d7e00000000,
103'h12eb277adf794e268000000000,
103'h0ec81845729f92bd72440802b9,
103'h0ca979b2c48aba385055fddd6a,
103'h0d2e92179252d27dc2bf693fe9,
103'h3e90e809defc4c308600000000,
103'h116c8c22ac2ade4818a0d6ed4a,
103'h12e7c2f8eabbc651f800000000,
103'h1aedb4077b285274a400001db6,
103'h33467793ce10156d8f00000000,
103'h2a9b8750a8fdc9750a00000000,
103'h0e1b75559b444108d80020804c,
103'h1f5729ac86dfc8598000000000,
103'h28bb307814fb3daf1a00000000,
103'h002f4cb13252675ba040da0669,
103'h00a1325f5b0d97d3b6d7651988,
103'h1a5759165a3ce484e8000002ba,
103'h3ced4826dade16e44400000000,
103'h337e74e676356ffa9f00000000,
103'h1b620901b322b8217afffffffd,
103'h1f5334f0a4a12d07f000000000,
103'h3e8145647f033609a200000000,
103'h388d6cbc9f566afa4600000000,
103'h28cf040f5cd7b05ec400000000,
103'h0b33538394651d1b6200004cd4,
103'h1138cfffbc34212abe82576a7f,
103'h15418285866774ae5200000000,
103'h38a0a00596a044ae0e00000000,
103'h36d76de46ae1c7339400000000,
103'h0a7358dea28267392a000001cd,
103'h194365039b59d51d9600000000,
103'h2f7ae5d6e4cd2dfc3800000000,
103'h1852ab583c1092ffd200000000,
103'h2e0c380d2a8b78d6b600000000,
103'h29482bfb44de242ef400000000,
103'h3addf506f2ea5c3c1e00000000,
103'h3240ec0eda3288376300000000,
103'h26b4761697107d3e5600000000,
103'h04b378f50851694d3000000000,
103'h2890a0026e05df63c600000000,
103'h3e58234bf2b95858ce00000000,
103'h2e522eccda49f85b3c00000000,
103'h365cb78c18a21ba73000000000,
103'h04b8a99888f44a740a00000001,
103'h031a7b08bf51020024117c0000,
103'h3235a4d1c309ab98ad00000000,
103'h3c9ac6f6052426a16b00000000,
103'h20a204c17659cb732c00000000,
103'h0c9d8d00f4f49269327ecfb4fb,
103'h36ea17409496972aa800000000,
103'h25404d18e234242b9c00000000,
103'h16baa992991e3b6c3200000000,
103'h3e8ed17f7d5e88851400000000,
103'h1c578bd592193217ac00000000,
103'h0eb6dd5652a803972a50008b01,
103'h234a5302aeff8f6cbc00000000,
103'h0efc041b3cb66cc30e5a020186,
103'h390c3db8de00bfc5bd00000000,
103'h3635a96e2cfcc3e0f800000000,
103'h050718baa6090199d600000001,
103'h02d81773dd3eab0804b02ee7b8,
103'h3a5f82f02145c3c2ab00000000,
103'h12e7ae32231ddb368600000000,
103'h176c9d551e7d5e26a600000000,
103'h00fa8e11f1650c58ca2fcd355d,
103'h06c729d6c6d1a9ade800000001,
103'h2cd9895e46cc37bfd800000000,
103'h3709c41c4c9361969e00000000,
103'h1eb75d00f96ceaf4e400000000,
103'h36ca023e7176af113000000000,
103'h14ae5129ce2e0c122800000000,
103'h395ed7d506f80e509900000000,
103'h28a2c016daa65f7a6800000000,
103'h1353934d9505374f6e00000000,
103'h2a7b15957ca7f7664800000000,
103'h12d0a3ef8efb8ab3dc00000000,
103'h011e409a3b76a0495a4a7071ca,
103'h0a123cbf4c474438e800000091,
103'h270b7033ce6584d32200000000,
103'h00ac9b0e9977c19270122e5084,
103'h2a49509d3e8331c63e00000000,
103'h0d5ca675412fccd4d6bff77aeb,
103'h3cb740862a791d721400000000,
103'h3a775f6a36d5c3e75400000000,
103'h10af3fe0b48d046d7e111db99b,
103'h266a521d6f0463d7b600000000,
103'h3b55312f00b3a3b86a00000000,
103'h3ab92db2a61df5d5d900000000,
103'h30f2ee1da0732704d800000000,
103'h1ab9b2f61a2c54b77e00000000,
103'h3284dba64b1f42d52100000000,
103'h0c03a80ee4d8f5cb3a6dfee7ff,
103'h0aa06a4d595dd171860a06a4d5,
103'h2ab05390a46179806a00000000,
103'h26ec918b6e01e3cdc200000000,
103'h2d48125b5ab2375e6600000000,
103'h177c88f6809ec8e9d600000000,
103'h1b0ed1032ce6db4530ffffff87,
103'h000292904363643bb0b2fb65f9,
103'h16f837eb1d72353edc00000000,
103'h06a014a45e74c7cf1e00000000,
103'h36e6ba47756cffba3c00000000,
103'h13143b2fbd0d145e9a00000000,
103'h32a52053b2f3cea60f00000000,
103'h2ea83ab6860809d5ca00000000,
103'h09201ce878ad2a297ec69b6083,
103'h1704fed4a75564e00400000000,
103'h22f6f51f6f7581c87c00000000,
103'h20dcba10457a809d2200000000,
103'h24ca88d6e77175bc9000000000,
103'h206581c7064e2fccd400000000,
103'h0255df972b18b8a3bc40000000,
103'h12bbbf2fca7e3a6ac200000000,
103'h269c1f658cd41a01ee00000000,
103'h22edf557de8fd931b800000000,
103'h268dfb17072bf8974600000000,
103'h1446b979e819edef2400000000,
103'h0c7db2478ea7e9062a7ffda3d7,
103'h1288c51722eea2801400000000,
103'h3923b118706c54c7a300000000,
103'h22ea95b102f519dec600000000,
103'h36cb6838bb18caf73600000000,
103'h1b5423c69e0360a838fffffffa,
103'h20cb81d494cec8e0f400000000,
103'h16af34aa2f22eca79200000000,
103'h0e88015e8eee6e7c2644002e03,
103'h0279990a249da3265664289000,
103'h156e915df425a484e400000000,
103'h3c325292b69f3d8f0b00000000,
103'h1319006f0d0dceecfe00000000,
103'h36ee1cc78840217fb400000000,
103'h0160dc465a5921eec0dcff1a8d,
103'h3ef9404a10473eb64900000000,
103'h3530e1dcd2a81afca200000000,
103'h3476525c90a15b46b400000000,
103'h3efbe45c04d23d238700000000,
103'h20da984a3a488f801600000000,
103'h15008aeeb94473dc1c00000000,
103'h1ace988fd91f0c2656000ce988,
103'h333e0177af1f97150f00000000,
103'h0e7fa78308ee2fa4e63713c000,
103'h2409dd0e7a2c311c9400000000,
103'h32d8867608abd89f9f00000000,
103'h18c63c03ecb5b5ae1800000000,
103'h2ed388a6de8e3c242200000000,
103'h0ccf04eeb85478280e6fbe775f,
103'h24f6b253272800ceee00000000,
103'h06ca385732f705bda600000001,
103'h1653740956edb810cc00000000,
103'h056aebdf9eb7f067fe00000001,
103'h2ad6dbddf40b64715400000000,
103'h376accab38765050f200000000,
103'h34f5c336224d2c2ee600000000,
103'h096e71d1d8b7f8da1eecc485e3,
103'h3c9f10d58cadbc104100000000,
103'h22db144a941c2de21800000000,
103'h028d681090bb3eb7a421200000,
103'h028ce805749653023a40000000,
103'h1d4460d47623bb12ca00000000,
103'h00a995b3b8b0a3183ead1c65fb,
103'h3a2af87514f503ecb400000000,
103'h076799ee169e99a06e00000000,
103'h043a8e6950c992158200000001,
103'h3a313df756312c039900000000,
103'h28d8909d9d6bba6cea00000000,
103'h2b74e730969cf8644000000000,
103'h04afd763fe758901dc00000000,
103'h2eb459ace8ea70327200000000,
103'h2eea07f96c9a47967000000000,
103'h0c8b70b2db4ea1435ae7f8f9ed,
103'h3ec9d1d08a38a93cc700000000,
103'h317dbbf016c419efa200000000,
103'h0a1c1642148debc02c00000038,
103'h1054b82a850ba7b042a4883d21,
103'h32dbfb564e27bdf25700000000,
103'h1e9be7bee17c761cdc00000000,
103'h201fee17125871732a00000000,
103'h3931e02f72f459320b00000000,
103'h144f79f8131447491e00000000,
103'h3e94d1b30b4627789000000000,
103'h0a569f8ade95a170a2000015a7,
103'h2970ded5df2a7323ae00000000,
103'h397f7752e88112ae8d00000000,
103'h1aa2571910f1f1846a00000289,
103'h090b5e57c87168d752bd1b404d,
103'h160a07072213bff06200000000,
103'h013322da2c1f1e482aa920912b,
103'h14dd515bc329254f4e00000000,
103'h36797161c35c48297a00000000,
103'h2286fa3f173999853c00000000,
103'h30a8430cceb30ae6fe00000000,
103'h2ae8aa22b13a05261600000000,
103'h27523687e0e24832e400000000,
103'h25180b168acaf2559400000000,
103'h3b17792a711d28dd7400000000,
103'h1ec9f225553533f3fe00000000,
103'h32b67046514cad1e6f00000000,
103'h2685369a2e169f43c200000000,
103'h251eef43a2cd0f8a1200000000,
103'h12d5d0ca895246244200000000,
103'h16c1e6456f713567e400000000,
103'h28faa8dec04706326c00000000,
103'h2a4a0abbd608ec77da00000000,
103'h0f667c23010395569c810a0100,
103'h3cd533ae6a4da0127200000000,
103'h16b520a1bab41c357200000000,
103'h32dc13c776894fe3df00000000,
103'h260bf3650d3e70859800000000,
103'h193f6859411a844d0e00000000,
103'h36c07d5fe62677b21a00000000,
103'h0ef5ae9bfe65e00b5a32d005ad,
103'h1cb42fbbf6265d6b4000000000,
103'h38b12161851c0c074000000000,
103'h12c8975422d03bc33600000000,
103'h150684f8da815d24ba00000000,
103'h14aa52a8ec49f478dc00000000,
103'h0a747dc440507971b600000007,
103'h045ab4e6d4facc1aa400000001,
103'h221127cc9e6f49dee400000000,
103'h1948f7d724c9fec5ba00000000,
103'h3ccabc5a86db26925900000000,
103'h229cfa4f9e241e697c00000000,
103'h1d6a045f5ceedac40200000000,
103'h34a6584dfe8bd513a200000000,
103'h32acab025af5d972ff00000000,
103'h348e24490e9c31c0fc00000000,
103'h1693bbf94148dcc35600000000,
103'h14882e6d76d7010c6400000000,
103'h100875f54d6abd05a64edc77d3,
103'h277e96f022f2eb731c00000000,
103'h0c90e9abf2fb6168687df4f5fd,
103'h32ec192b1a79f8588b00000000,
103'h0f1e49b6a70ae2047e85200213,
103'h36bb3747d8f6fb2f9800000000,
103'h034b104c271544e63e80000000,
103'h00d64ab8dcd07c2e16d3637379,
103'h18db7d7e1f1b8c7a3c00000000,
103'h16eb9247def1d7331800000000,
103'h2cf2a24136cd54b13800000000,
103'h280ef720ccb8e6f91600000000,
103'h00fbc82e78ab893a4ed3a8b463,
103'h380425b660ba805b1b00000000,
103'h10fe5a7162b64889942408f3e7,
103'h1ec5e3dd9aba6e3ff400000000,
103'h38465442eab8c8b15700000000,
103'h0c724de2897eac8ef2bf76f77d,
103'h0358c7dd42c500d1dcfba84000,
103'h18f58a618f374eb46600000000,
103'h0a4cbb25d0901691a800000265,
103'h295cb49b6a85a0f33600000000,
103'h0eeb5a9ff4d25c1908612c0c80,
103'h363f01765d2f10b47200000000,
103'h2cc9f7012a1a6b546600000000,
103'h34e5031da1596ccac400000000,
103'h2685b02d4e2363cbee00000000,
103'h0ef8b956030866e99004102000,
103'h129ad3332a8e1716de00000000,
103'h01575864b886d06ce0ef1468cc,
103'h116d4a610a21a3a00aa5d36080,
103'h2ea6a0294a78fc04c200000000,
103'h10e85cdb1ce64665cc010b3aa8,
103'h1ab830a3ca8ce68f180005c185,
103'h1e0ed4d95b75436a3400000000,
103'h2a871caef62d740dfe00000000,
103'h03786089553c48e75a08954000,
103'h364feac97ec365965000000000,
103'h36b45b98c33bc61fa400000000,
103'h108e0fd2388bb0e922012f748b,
103'h20953819ae400c81e400000000,
103'h04d8a9487ece1c541e00000000,
103'h26df800d9e63546dcc00000000,
103'h0c221cf2633bfdb64c9dfefb37,
103'h2af06ac04a1b7dc3ea00000000,
103'h36fec510173d9ab64e00000000,
103'h02db3bb4012e057698dda00000,
103'h2e1b06c5b72cca86ae00000000,
103'h3c96cf8dbb08063aaf00000000,
103'h152e1619a8230d006400000000,
103'h0302f75be4b9dc8e1ed6f90000,
103'h3105de14b8e7f2a7c600000000,
103'h15358f543aeaea03aa00000000,
103'h356d46ce6af0c8186200000000,
103'h3ac80b48fe26576c9d00000000,
103'h26dcac51b2939e3b0600000000,
103'h08d940022f5ba98406c174c314,
103'h26c0bdb6543855d5b800000000,
103'h2c990382dc1195d7e600000000,
103'h3297a0bc02d2538e3b00000000,
103'h2d29dc30316b57111800000000,
103'h1217c1286202f7cd1a00000000,
103'h0e3dfbf64e2cd3fd4a1669fa25,
103'h2775cc9c23449525ae00000000,
103'h017ff0d03082911bfc0140f616,
103'h0cf56c1556f85db81e7ebedeaf,
103'h3a6ddf2796784e884e00000000,
103'h36132637226dba9da400000000,
103'h16fd026c5cdb99c53c00000000,
103'h25696fbd94eebffc5e00000000,
103'h0ace3ac6eaebc268bc00000001,
103'h06ab54588f5532265000000001,
103'h24f62887d9236ced3a00000000,
103'h201c967c5ecec145c800000000,
103'h3131c46d44c4e9cda200000000,
103'h2a32b4c6e4e1804a0000000000,
103'h3488d746d61344b74400000000,
103'h160266b40145f97e2a00000000,
103'h164ab766f4ced0c50000000000,
103'h1c57f1e78ad137790000000000,
103'h0746acb2231beedff600000000,
103'h0748ac33fe73e0c78000000000,
103'h0690a53404ba8d79a200000001,
103'h3ca76ef90a0339ada000000000,
103'h3e8f70371093dee1a400000000,
103'h209360550e3b4ddaae00000000,
103'h030b313a8ccabe11c085989d46,
103'h263d8f99ad5e1e66ce00000000,
103'h167327a66f694fa15a00000000,
103'h173c9e94d6a6df3b0600000000,
103'h2541635ded1a06e17600000000,
103'h3f10e638c356a5764c00000000,
103'h053e877a669808d43800000001,
103'h3ad5785d64a8ef0cfb00000000,
103'h0613487b68e776876000000001,
103'h3f6b1f7ae4bceee4c500000000,
103'h38199bf0aad037602d00000000,
103'h1960213aaa3b56db1000000000,
103'h1c4f9591a354f2cbbc00000000,
103'h0b26806ffcb514066600001268,
103'h1aba5a331804a9980805d2d198,
103'h161e6b56622b2a080400000000,
103'h3cbdd354bee5843b1f00000000,
103'h06b22e1ed403ef918000000000,
103'h0b5b9cef52c1c2e63e00000001,
103'h2909b557d973f1051400000000,
103'h2ae2f7c862cf8df46600000000,
103'h28a1be740cd9434c3e00000000,
103'h3d6474b136bc3b14a000000000,
103'h22e8edd49e5df988ac00000000,
103'h20e157fd1cc26e39e200000000,
103'h02a95019feab5c0e82a95019fe,
103'h2f4a8b83208cb40b9e00000000,
103'h12a80200e23604259c00000000,
103'h1463720750808fa8bc00000000,
103'h32e15047a22891a99f00000000,
103'h0e0a8a96768c03b0f004014838,
103'h0cc078f0e86d53f89276bdfc7d,
103'h2aac6b70f977de8f0a00000000,
103'h1b18ed99c438577ff2ffffffc6,
103'h2eae016c2ee4c2f0ea00000000,
103'h38cf18ef8afdb08aaf00000000,
103'h2b5d846b78abb1f6de00000000,
103'h1763ce76717acae66800000000,
103'h04a270015ad84f51e000000001,
103'h22c5d47d313c1dc85000000000,
103'h0ae6e983b6de8dc9aa0000039b,
103'h2ab3b08118a46246dc00000000,
103'h3afb4264e48b4bca9300000000,
103'h261b239a8e3efc4baa00000000,
103'h037722988a3a3eb08ec8a62280,
103'h14b1af603155624b1e00000000,
103'h3e909e6eb2cc84e3a800000000,
103'h0efad947c77e3443d83d0821e0,
103'h2ca4106c850ed2b28a00000000,
103'h14878641d309abfa5000000000,
103'h2cc05e623eadbc66d400000000,
103'h36c5bb66533542a8a800000000,
103'h06494cae3ef5a10ae600000001,
103'h1adbb0a8b4bb5c713a00000003,
103'h0277c09d7a04a91f78d0000000,
103'h2ac18cf916e059c82e00000000,
103'h24409bfd58581a65a800000000,
103'h1cb54c0c8219a75ebe00000000,
103'h0ae5588ce75a435c1800072ac4,
103'h351a0e2cc40f8f689a00000000,
103'h322f1d94cef4e7f58300000000,
103'h0a9c4762830ef6224609c47628,
103'h2723188ef63e13b71400000000,
103'h28042d1780da5b199800000000,
103'h2ef4d108a6fd73a88e00000000,
103'h02da5cef4e01a0c00e973bd380,
103'h1acedef83cf671c8b60000000c,
103'h290174b840d0ceb80400000000,
103'h380e6591da9fadb04300000000,
103'h2f18ca1404a122688200000000,
103'h3324cf563caf87fa5d00000000,
103'h352746612ac8520e6000000000,
103'h36fa8c241ced21649c00000000,
103'h156d7f97521467c5c600000000,
103'h34819573090ef3e9e400000000,
103'h124533491d7c73813600000000,
103'h18d1232d92fe08f43e00000000,
103'h3d4a3476a5433c3d5c00000000,
103'h32d7ad857d145f6aef00000000,
103'h33741a7e3b5e93e19300000000,
103'h0e8cfaf82c3641670e02203006,
103'h3ca3e4665eaa5be54900000000,
103'h0efe0a11ed3756dd761b0108b2,
103'h1c6c8f2868db3b43d400000000,
103'h2639a82076d94555c200000000,
103'h1d3d027f9445d47e2a00000000,
103'h30eab8c3fb7f7c9ea200000000,
103'h32cfc5e5d6bc7f1e3700000000,
103'h1e900e4b86a737e23000000000,
103'h01299c06fb76fdc806504ce780,
103'h3708fe4098070c138c00000000,
103'h2767dd18d830a81a8600000000,
103'h2c833b0f4e39a65b1e00000000,
103'h3945d0e7f4a18373f700000000,
103'h017f6488a024be8344d21185f2,
103'h1ec0043cd86a8f6b3800000000,
103'h16314c0b98e9f3f3d800000000,
103'h1adc3a3578a9f830b200000037,
103'h1528abd34edb443c4a00000000,
103'h2c99dbf468b77e71c200000000,
103'h1e759b80bce02a451000000000,
103'h2b3b4f00eb7a06397a00000000,
103'h2caafab1c8efa1ba3600000000,
103'h3ef5ea9ef22af0bb2100000000,
103'h38f858fde0d5eb6cea00000000,
103'h2edaf1a1decbd60bdc00000000,
103'h1137907f56c42f09bc39b0bacd,
103'h3a83d117049f20ab9a00000000,
103'h16fb0269d4d6b12af000000000,
103'h14481f298f5a8241f600000000,
103'h2f6111f5265584abca00000000,
103'h213e33ca7a9da3d55a00000000,
103'h16ba764b68feb5ca8000000000,
103'h200d69f7493ce994fa00000000,
103'h3abadfe51ef75fe06200000000,
103'h3abdda7ec104c9d7ad00000000,
103'h345e78edbabfa9bcca00000000,
103'h18fdcd27367d843b8a00000000,
103'h04da0af5aadbfd294600000001,
103'h0eada8a482d9ca507c44c40000,
103'h1a86102b06b3d5462600000861,
103'h211e216e57617deaaa00000000,
103'h1d33b6ed30e78e15b000000000,
103'h032549955005af840695265540,
103'h2cf0a68dec3966713600000000,
103'h1e6fd8ccae5eb0068600000000,
103'h255088f61c4f56947200000000,
103'h1d18c7353abf2f612200000000,
103'h22e6b4f85f0fb8573e00000000,
103'h16ee092cbb287f8c7800000000,
103'h39540d679e0f3484d700000000,
103'h37096836f4fd3db19200000000,
103'h2f7df2676d514b193000000000,
103'h050234ef235ab3502400000001,
103'h16aef70350d8a5b79000000000,
103'h066aed9c54dadaa6b200000001,
103'h2b2421e6ec89d1aa0200000000,
103'h3a2ea14ab2f4bf465600000000,
103'h2c93d3fe9e18e12d4200000000,
103'h2ed1ac6a19478277f600000000,
103'h06ea5f7c46db56769400000000,
103'h088ce43874ad02e0ac10f36c6c,
103'h3e24283afa97625cf200000000,
103'h12d44d6ac52446956800000000,
103'h00cbf51282486ed0628a31f172,
103'h329ef330d61cbc3b2700000000,
103'h1b1ef42fd6e8b14daafffffc7b,
103'h3e36578bc887a47e8000000000,
103'h2572017d24a698ae5600000000,
103'h0ef61a3ee2dcf03a1e6a081d01,
103'h0e96ef3bc64ef1b742037099a1,
103'h2520758656450bf62400000000,
103'h0431a04f64dbfb31ec00000001,
103'h06e963c6cafc70b84200000001,
103'h2d7e17784e2e1107a600000000,
103'h1861bce1141774ce7000000000,
103'h1a8a6e4000958c46be00000000,
103'h008f1ad0d8f74927d4c331fc56,
103'h32903819f281b767d500000000,
103'h30bf666ab510d238ae00000000,
103'h05060989e6a10a52a000000001,
103'h1ae238efd66070bd54001c471d,
103'h08b5b17d9c667a473a69e59d53,
103'h290ae1733748b3371200000000,
103'h3f70e3a17efe64b4af00000000,
103'h3877f02267094627e400000000,
103'h0adf6d60a57a29c962000037db,
103'h38ad64e61ef219ebc900000000,
103'h1cc40fa2a8d1874c6e00000000,
103'h3ed91f13e37eec328c00000000,
103'h08f774acfe42fbd5345ac7bce5,
103'h368ff40f7e1c1ae91600000000,
103'h031a8d5dc7138f961635771800,
103'h3776adf87ca383a59400000000,
103'h0f51bac5bebe11035a0808008d,
103'h246fc3683534befbd600000000,
103'h38a9e6f3c28679c19400000000,
103'h12f79a1566f63d29c800000000,
103'h28e8d0dc9ea0241d8c00000000,
103'h3c9818a73097be32f200000000,
103'h047c1f6d98808f0f9200000001,
103'h10e69ff59418a7b6c266fc1f69,
103'h05475da75a94c7245c00000001,
103'h16483f76aa7b6719f000000000,
103'h18e0df78eec2c4c14a00000000,
103'h34fa0e8ac50b0437f600000000,
103'h272be5535eebe3b0e400000000,
103'h30f2834052e5f23baa00000000,
103'h263488473911d78f0800000000,
103'h0d39520f6a045acf5a9ead67bd,
103'h3649200f9138e3169400000000,
103'h3e44d1c09d723525fe00000000,
103'h182675ad52bb55358e00000000,
103'h2c19f129110026f62c00000000,
103'h2b11c7742a269ca37e00000000,
103'h3a4280d5d7408dcc9100000000,
103'h26e56f5d83525540ba00000000,
103'h2543b31abc94d6169000000000,
103'h34a21dce227a45741200000000,
103'h2e27252506bdf88ece00000000,
103'h00ecba487c60165cf0a66852b6,
103'h1204a4acaa873b81f800000000,
103'h22b165276b73f5ca7400000000,
103'h12d86b163e789a771e00000000,
103'h0abd6993e129ff9e8a02f5a64f,
103'h3e027e6e73026ab4c800000000,
103'h1ecececafebfd448a800000000,
103'h280f14f1fcc252b71a00000000,
103'h30c7f5901a9121821800000000,
103'h18aad5ccc2a036741600000000,
103'h329020be32682c043100000000,
103'h0c353ff84b1301d0f49b9ffc7f,
103'h229cb1e97ea3228f2600000000,
103'h1295455ccad862877200000000,
103'h072e0f442d751470f000000001,
103'h2e2f052fbf0a59cdba00000000,
103'h2142fcec47386911e600000000,
103'h10fa1737f4676e41a449547b28,
103'h0a89940b14aa6b2dea00000226,
103'h308e254f24a48265de00000000,
103'h149d1060ee2e1670f200000000,
103'h00e464849ebc3bc016d050225a,
103'h1e9326e9f2594c210400000000,
103'h12ec547d323db0a5a200000000,
103'h28ea047652d0d78f9600000000,
103'h2f15cae064bd2c0cc800000000,
103'h10fdcd0a8ca730831a2b4e43b9,
103'h263f1b55babcfb637e00000000,
103'h30be1a468cbac86e0c00000000,
103'h0a0df0c6f2f9e3c3c600df0c6f,
103'h0a1af35422b7fe0a520006bcd5,
103'h16cf26646ec5eed14600000000,
103'h1d4054d838e0e2256800000000,
103'h316c4bba0eb00889d600000000,
103'h3692265faaf05d620e00000000,
103'h1e6fff0f9a5ca91c1c00000000,
103'h3613c690d0eecf7bc800000000,
103'h04987037705ece8b6200000000,
103'h22cd2267e772951c3400000000,
103'h2af231fa6b0b0553a400000000,
103'h0c73eaa90cd827bb8a7df7ddc7,
103'h00e472d376ca59b5f4d76644b5,
103'h24b3c989453e445f0200000000,
103'h2ef5b55b4422b7327800000000,
103'h2542a680ead680bbbc00000000,
103'h2667bf6218cc36170200000000,
103'h1e5731f93d0edc97ec00000000,
103'h1c84e8ef62769bfa0400000000,
103'h1ed5571802cdcdf34200000000,
103'h0afc45fc5e52b6e2a400001f88,
103'h0eef6af7bc280dfaa614047952,
103'h10f16c8b062453f704668c4a01,
103'h366a0a185413beeec000000000,
103'h1cb07598e6052b79c600000000,
103'h234997fc1d6f35921c00000000,
103'h220ac859f91fab2b0200000000,
103'h2af04caedb6943271e00000000,
103'h06e98ff27e740b811600000000,
103'h08e7feafe964582ff2c1d3400d,
103'h2755a2ff6f4de8227000000000,
103'h3ce2f279f735e6d25900000000,
103'h2ed9851b9c8b89d1c600000000,
103'h1e44233e596e7c4bbc00000000,
103'h37131991094801675800000000,
103'h3c2ff806268c24a5b100000000,
103'h3882bd4d9e9f3e36b900000000,
103'h10610c66dacf363ce0c8eb14fd,
103'h02add7cbd551f38a7e00000000,
103'h3a42a49824b2fff15800000000,
103'h1a63960a2660d7bd2c000000c7,
103'h1923c5b2e2a37c555200000000,
103'h32b32b987c07125f7900000000,
103'h1e948508962ad8125a00000000,
103'h3128de6a08de03aad800000000,
103'h2a1e0f88a77288b36e00000000,
103'h04b6bcfc989b671d7600000000,
103'h1d567cd002b976a61c00000000,
103'h0a2114b5c67033a2b400000004,
103'h00c9b04664c6b072b6c8305c8d,
103'h1ee4d48a6ee7c5287e00000000,
103'h129b5febf0b1756ee200000000,
103'h0b0b61f38e9649f9500085b0f9,
103'h08eb979de031a9e5406d1f3c50,
103'h2a927dbaea3d0bd8ce00000000,
103'h3a2129007328a376b100000000,
103'h3c6149b4dcbb21319b00000000,
103'h0b37b46298dc4a320e0137b462,
103'h3b3fc8f5943d93e6ea00000000,
103'h1684e9615e7548498200000000,
103'h24f2ad43dab5113f1600000000,
103'h0f1b9257f139faa0768cc90038,
103'h1320c19e152ca7e45000000000,
103'h286384cb23483a3c4000000000,
103'h1e1b9041b568fbda5400000000,
103'h2e88acf75ecc80a57600000000,
103'h2e2fc44d7ce810e72c00000000,
103'h03038387ed70bdde8a38387ec0,
103'h3a1f7cfe9aa0822c0600000000,
103'h26a4724f9ea405b3f200000000,
103'h30f5e84618c382b28e00000000,
103'h372f6f23bf67f5022c00000000,
103'h2ad9b3dfef5ddd484400000000,
103'h38247ac8248d4c6c0300000000,
103'h241347644f67004bf000000000,
103'h28c596b3068b7b141400000000,
103'h2adfdb03ea9ec2786400000000,
103'h1a57fc9d1264592b6a0000015f,
103'h2e5d6aa23d44342f5600000000,
103'h12c9d8f3569c30cc6800000000,
103'h3ec1c25886f99b6ea600000000,
103'h14586e3618c37461fc00000000,
103'h3c53733f168536ba8300000000,
103'h2292ac776adda4f09c00000000,
103'h216e167c2831182fb200000000,
103'h22431bef8ac3c4a71e00000000,
103'h3edb95c4eb31db234600000000,
103'h32f94654ce74f712d100000000,
103'h10f49bd54d508cd7bcd2077ec8,
103'h162109857f49d32c8a00000000,
103'h26113bdcce3e6f01d600000000,
103'h22334957655f78875600000000,
103'h2cca4de4cc70b4642400000000,
103'h04b1df49eea3fdbb8a00000000,
103'h1ae343db9d6e4ba056000e343d,
103'h3f53176f20202aea4500000000,
103'h09226389fa036ec5e09086a60d,
103'h1e626408f85686350000000000,
103'h254662438278e9befa00000000,
103'h0498ac1e60db4dc7f400000001,
103'h060b20e38521b00b7600000001,
103'h0081046e8aba5c29d69db04c30,
103'h354d6e2e90c57d0d5c00000000,
103'h2a92c1ad9146817be600000000,
103'h02b362f48693efaa7618000000,
103'h1ef5b446f026b1580600000000,
103'h04f261c332da144c8c00000000,
103'h3ab48c4cd0cfc8937e00000000,
103'h00bd385254c22a56b0bfb15482,
103'h0e59d4024f76b6a382284a0101,
103'h0d1d210a5033eef5d69ff7ffeb,
103'h3cba825ede8dc2f82600000000,
103'h3f27ac46eaaae4027700000000,
103'h16570085a76566615400000000,
103'h3cfd0b67e68d12a83e00000000,
103'h32d7053ffce4132de500000000,
103'h073ec21038e11e95ca00000000
};

endmodule
