module uart_tx_sb_ctrl();


endmodule
