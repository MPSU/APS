//////////////////////////////////////////////////////////////////////////////////
// Company: MIET
// Engineer: Nikita Bulavin

// Module Name:    tb_fulladder32
// Project Name:   RISCV_practicum
// Target Devices: Nexys A7-100T
// Description: tb for 32-bit fulladder
//////////////////////////////////////////////////////////////////////////////////

module tb_fulladder32();
    timeunit      1ns;
    timeprecision 1ps;

    parameter TIME_OPERATION  = 100;
    parameter TEST_VALUES = 3000;

    wire [31:0] tb_a_i;
    wire [31:0] tb_b_i;
    wire        tb_carry_i;
    wire        tb_carry_o;
    wire [31:0] tb_sum_o;

    fulladder32 DUT (
        .a_i(tb_a_i),
        .b_i(tb_b_i),
        .sum_o(tb_sum_o),
        .carry_i(tb_carry_i),
        .carry_o(tb_carry_o)
    );

    integer     i, err_count = 0;
    reg [97:0] running_line;
    reg [98*3000:0] line_dump;
    wire [31:0] sum_dump;
    wire        carry_o_dump;

    assign tb_a_i = running_line[97:66];
    assign tb_b_i = running_line[65:34];
    assign tb_carry_i = running_line[33];
    assign sum_dump = running_line[31:0];
    assign carry_o_dump = running_line[32];

    initial begin
        $timeformat(-9, 2, " ns", 0);

        #1; // wait initial line_dump

        $display("START simulation of 32-bit fulladder.");
        $display("You should run simmulation until the message 'FINISH simulation' appears in the log.");
        $display("If you don't see the message then click the button 'Run All'");
        for ( i = 0; i < TEST_VALUES; i = i + 1 ) begin
            bit fail;
            fail = 1'b0;
            running_line = line_dump[i*98+:98];
            #TIME_OPERATION;
            if (tb_carry_o !== carry_o_dump) begin
                $write("ERROR! time == %t. ", $realtime, "Carry mismatch. Received: carry = %b, but Expected: carry = %b. ",
                    tb_carry_o, carry_o_dump);
                fail = 1'b1;
            end
            if (tb_sum_o !== sum_dump) begin
                if (!fail) $write("ERROR! time == %t. ", $realtime);
                $write("Sum mismatch. Received: sum = 0x%x, but Expected: sum = 0x%x. ",
                    tb_sum_o, sum_dump);
                fail = 1'b1;
            end

            if (fail) begin
                $display("It should be: 0x%x + 0x%x + %d = {sum: 0x%x, carry: %d}. ",
                tb_a_i, tb_b_i, tb_carry_i, sum_dump, carry_o_dump);
                ++err_count;
            end
        end
        $display("Number of errors: %d", err_count);
        if( !err_count )  $display("\nfulladder32 SUCCESS!!!\n");
        $display("FINISH simulation, time == %t", $realtime);
        $finish();
    end
initial line_dump = {
98'h04854d49302257a06d29e93a6,
98'h2c7c1598c1ae5ec36b8a9d171,
98'h2cb0a119624dd484b3bf9d678,
98'h01b5f3434ec8fc5da41fbbe84,
98'h1db515fb518b7de32bd024f7a,
98'h38cdc931b8bde1315c62ea98b,
98'h1cabfdf96ef49c9dd2e826a5c,
98'h11fb36e3de4c1a7c8c11d4581,
98'h3d001eba38b293b15d6cac9ad,
98'h37a38a2f65aad60b7753980eb,
98'h2c7bd898c15ce1c28b762e96d,
98'h04190848155e116aa65dc66cb,
98'h32c80fa5a260ee04f54a3f6aa,
98'h2a69f594cd67f75aedf47b3bf,
98'h2045d280b5d58fabb586d88b1,
98'h39f15cb3c4611248cf949bbf2,
98'h395cc2b2a78c530f183a45706,
98'h114b986288312cd0465f314cb,
98'h0f083cde312284a2700ab0602,
98'h16c0996d98d2fe718be4e5f7c,
98'h379d40af0543f74aaf384dfe7,
98'h2e25ef9c50bc90616fb89fff7,
98'h2773180ec7418cce8bad29375,
98'h02aa92c55e3666fc68383e707,
98'h0c48c1d8898d7ed32575902af,
98'h11ee6863df1b6a7e2c4274b88,
98'h33f115a7eb9f651737e41eafc,
98'h11378de2692b8c924e98c69d2,
98'h3affb035ea31ff14594c6bd28,
98'h01875fc3384b33b08e74a4dce,
98'h2ee0969dc7bcbb4f4da7547b4,
98'h2fc1401f8db9605b6f5ea81ec,
98'h03f4a3c7fa7afdb4ef9be85f3,
98'h2f05221e0b769656ee9eee1d4,
98'h27fcab8fc5432bca8b4ff5d69,
98'h30cfce21b1c6832398a594514,
98'h1f4d667ea4df6f09b10b35621,
98'h3462ed28e5e66a0bf69255cd3,
98'h2bf61597c88a43512d20163a4,
98'h3966cdb2fcc246b99d8a451b1,
98'h0533f04a7da0b8bb50b52a416,
98'h2ca7ed9976a2b8ad78d2a991b,
98'h0f3c465e488c7fd105f2318bd,
98'h054242ca957dab6ac6affb8d5,
98'h1b976b773357af26b3bbc6a77,
98'h387c40b0cac3bb5590cfff019,
98'h2cf65d99e14c4d029390aaa71,
98'h2703a28e0f3461de4d8e011b1,
98'h129d2fe512719764c943b1d27,
98'h2b2df2965b72da76f1a833435,
98'h1b2c2df66da9099b52354de46,
98'h194ed27296c5cb6dac0527781,
98'h28c1c691809d26c12a57bb54b,
98'h0d2601da769baead10f06c21d,
98'h051f364a25a4010b6ab0cdd56,
98'h25d7270ba11df90211bd48036,
98'h3fa9e9bf452781ca51345ae26,
98'h10cd59e1bb4d0236b30697061,
98'h0cd3a9d9ae15711c2eba46bd7,
98'h175c666e8bceacd788cac4d18,
98'h1aa3817563493d86af7b2fbf0,
98'h06e1d84dd2c9cde5866ae98cd,
98'h04c967c9b6d186adaee6bb9dd,
98'h1b97c3f710d855e18b1c06762,
98'h0fd6a6dfbb636036f2ce81c5a,
98'h0f3b4ade7f4a393eb3a161074,
98'h02e50245f43d5e284dc8981b8,
98'h2a18e5941ea3167d722eff046,
98'h2526a28a582c5d706f54bffeb,
98'h33006d26096c9ed2ef1b42fe4,
98'h3d88b9bb315405a29bb72fd76,
98'h3512e02a1527bf6a728ea7e52,
98'h01c2ee43bccd19b9afa401ff5,
98'h054bed4a8556874aa2a89d255,
98'h13dd7fe7a71b798e2ebe3e5d7,
98'h191938f21948d172ac9882993,
98'h0d68325af8edebb1d19587832,
98'h1741676e9885aaf12bf1c497f,
98'h124bf4e4b689a6ad323566e47,
98'h30cce4219f5b7d7e940a18680,
98'h0651484cb7b397af4f8137fef,
98'h3c9269391950f3f2b578d74af,
98'h34256a2851d96a63b17fb5230,
98'h21794782fde0a43bf7d67aefb,
98'h06d8394daeac521d6d6122dac,
98'h0d736fdad11979e207a33a6f3,
98'h137ce066d24f916489731c72d,
98'h25a1380b496dd7d2cbc3c3f78,
98'h23c73d8781acc143495cffb2b,
98'h0300e7461a2b86f4474b1b8e9,
98'h28300910676fd90ed3e7f887c,
98'h0a7bfa54eac65895ad5094baa,
98'h3c59beb8a09cf881373dadce7,
98'h3b142d36024f93448f58f01ea,
98'h2720448e7ca1edb978f08c91f,
98'h056243cad0241760456196cac,
98'h04ed5549d4357e686648b4ec9,
98'h20888e810b0b48d60ae4f5d5c,
98'h029ba4c522466d04893884726,
98'h362b38ac4ab0b5557036fb807,
98'h0562cacadeac46fd6903c4721,
98'h24f04889d0927fe12d60b21ac,
98'h3cf5e9b9f73be42e7d0c737a1,
98'h1b796ef6d92e83f26d29fcba5,
98'h342f17a84551b74a8e6033bcb,
98'h28b9881150684160ce48725c8,
98'h2e51851cbfd3cf3f9b8955170,
98'h2df7ea9bd0d183618fb25b7f5,
98'h071c65ce081da45003ce82878,
98'h1ec36a7db8afc6b155dccc4bb,
98'h0e9897dd07379c4e45740d0ad,
98'h078721cf054864ca8333e1a66,
98'h02bb0d457c2c53b86fb9d83f7,
98'h2862fb90d92d78f250641d20c,
98'h04a5f2c9583da7706738e68e7,
98'h2b59f89680f589c1cb13e0961,
98'h018297432e2b799c6beb8437e,
98'h16d8396dbef7f0bdd5740a8ad,
98'h2b9e16170aae3dd54d9314fb1,
98'h3402c4a80e58025c9096b1c12,
98'h1ba2bd7761b73c036f567e5eb,
98'h2f33109e73d8f6a7b8c301d18,
98'h2f78349ed1f89ce3f05c3460b,
98'h1c704a78c3a490c7680536d01,
98'h088467d132a72f254ecae5bd9,
98'h3da85e3b4a5e85549201b8e3f,
98'h11b72de36a57f1148f03c7bdf,
98'h08dabf51b18ea4a30e9a58fd2,
98'h02fab045cd4b585a841182281,
98'h3556ef2a8f9bc3df113cacc26,
98'h1752936eb1685822d22ebae45,
98'h24a0c789464160cc8ab88a157,
98'h2923df1262992c0532ef42c5e,
98'h097c80d2eb9a0c172d45a33a8,
98'h10cfa5e1a72bde8e4dfee11bf,
98'h1a1479742588940b0fe7435fc,
98'h00fa6dc1ed48901aab90bf772,
98'h1d1abffa2979e792f1a529e34,
98'h1d8a56fb047f8148c8827610f,
98'h193859726729c10e701886a03,
98'h3a9605350ce0d959f1ddb7a3c,
98'h160c496c10440e60a99415f33,
98'h3b2e46b644002dc80fcb9d1f9,
98'h126c5be4dc6d1878cbb65d176,
98'h391c7e322bb5cb97593492725,
98'h1089aa61256a6a0aed7d051b0,
98'h225fc704aa5fc014b32fe1c65,
98'h3a0ae5b42dd67a9bb9f85813f,
98'h1b62e1f6d4d49de9ac0ddff82,
98'h201e5f0021f91303f085dc810,
98'h2194d8830b2a06566b2fb7b66,
98'h19f5cd73d20e79642b0111b60,
98'h2d3e691a4ee0f35dcf07d71e0,
98'h3b0dd63613775366d3a14a673,
98'h171e2c6e36f9bcadd385fa46f,
98'h2613568c0efb54dded43aada8,
98'h1a857d7500e1e1c1c6d9d7cdb,
98'h1d286b7a5178a2e2eba843975,
98'h1b6022f6f01d90a012df6ce5b,
98'h38bb36b16609fe8c37b14d4f6,
98'h2cc0b69995feee6bf0afe9416,
98'h1f106bfe20ddab01affb85bff,
98'h1c3bcdf872ad1f2553ba3b476,
98'h0c1393583ca717b9522eaac45,
98'h0c8bdf59052d0dca646e3b48e,
98'h2eef149dcdc5455baf2d167e6,
98'h1aa7ee754d0df55a09ed78f3d,
98'h355e002a81e7f0c3edd17c3ba,
98'h2fa6ef1f51cba563905ca520b,
98'h0799934f352d79aa6f31c33e6,
98'h2b79f416f5e88f2bd858a0d0a,
98'h1734836e42638b44e66603acd,
98'h0cb710594a3189d465ba268b7,
98'h332604266744820eb69aa18d4,
98'h0c5f01d8bc8d5ab9123b17246,
98'h2fb6911f4b3b97d66ebc8a3d7,
98'h1db79afb792a003275b866cb7,
98'h15f0746bfb69c736f4568ee8b,
98'h0e04e7dc20c9b5018bb3a7376,
98'h17a60f6f6d55779a913ee1c27,
98'h2a1b17942f61bd1ef65f352cc,
98'h2f0fe11e1edee27d937bb0e6e,
98'h047326c8cf2ceade44e80469c,
98'h377451aee1c33b83b64de34ca,
98'h019c40c339c3e6338ed809bda,
98'h2b3b371657289bee7098f4c13,
98'h1e93effd2ebd389d53544a269,
98'h273f1e8e405ca4c0a9e6f0d3c,
98'h00befe4149c710d382a183c53,
98'h171e546e211fec822e0f903c1,
98'h35ed23abdd1ccc7a14c27c097,
98'h1ebdaafd69882413321173c42,
98'h2801699004aa40c96b2aea966,
98'h2e1f041c05b2fe4b6cf48099e,
98'h1789546f261ec20c0f6a059ec,
98'h0a1d9a543433daa86f945d3f2,
98'h3ebccbbd5ea1ebfd7757adeeb,
98'h329204a52d56299a97fa0b8fe,
98'h3710c22e33cc27279ab73a556,
98'h08d002d1a0fe9901ea73a6f4e,
98'h2ab69d1556f4f6edf06ae500d,
98'h2c600298eb24f81655e13eabc,
98'h2d125d9a23d8f907943ad5a86,
98'h0b4669568390e14723b5d2a77,
98'h156187eada09b6742bdacf97c,
98'h1b1a9b7628b3221170f36f61e,
98'h117cc8e2df89247f0c417b587,
98'h349fc2a90325e3466df1697be,
98'h27ce638fbe62f03cd98c54f31,
98'h18815af10b8d90d70903baf20,
98'h33475426830586462d93369b3,
98'h1545746a834480c6a6227d4c5,
98'h164d3a6c818cd8c325f684cbf,
98'h1876bf70dd6b5cfacd78871ae,
98'h1e4b00fc9120eb626bdafb17c,
98'h037852c6f5a84a2b4e48273c8,
98'h24be448959fa15f3efae169f5,
98'h23653486f00ecfa034dd0109c,
98'h104b7f60a08d10812c3623f87,
98'h06cda2cd865a80cca34a08e69,
98'h3c92ebb922d0bb0597d8e9afa,
98'h1814197025d6620b8f7a9edee,
98'h2e30309c5f7fa3fed36bf526c,
98'h3b9c1a3702fb15c5efa5cbff4,
98'h1d7ec87ad6a74eed6d0985da1,
98'h31ecb8a3f7fdbdafda7a9d94e,
98'h3a6d26b4fac740b59d4d19da9,
98'h0358dd468e39a9dc6464a1c8c,
98'h21d8a383be31c53c78029a300,
98'h00af50c1438ebac7010f82e21,
98'h3d9c223b2550758ab8bb25f17,
98'h06e4814de07e8d80c9d8c3b3a,
98'h3fab773f67de838f99e27eb3b,
98'h2e980e1d1602626c11269c224,
98'h02459344ad1abf1a2bd81497b,
98'h3fc80bbf86c3c34db1a2f3c35,
98'h1f776afeed635f1af336b2867,
98'h21f40d83e291ed8511217ec23,
98'h34d99ba9ba9d89b53bddc957b,
98'h2d61f09ac09dfac10b7ffad6f,
98'h11a2d8637c3a9c3873775d26f,
98'h37265d2e7937c5b25c1788b82,
98'h28d90c91879d32cf2c1d8fd83,
98'h0b0315560e7595dcc65e2accb,
98'h1b9b48f7060ff0cc086ace70c,
98'h001cf940086083d0c21f5f443,
98'h342e66a84a7007d4cfa79b9f4,
98'h0bfbcf57f0efa4a1cf3adcfe6,
98'h05a6744b6e1d809c2cf0fd39e,
98'h2635ce0c624bf00492206f843,
98'h01b6dac342b344c5411a87e22,
98'h1298e3650a86e8d50747f30e8,
98'h02634544f878e1b0eeb709bd7,
98'h3b93b9b72f1e041e3aac6f755,
98'h2bfb4997c47016c8ec1ad8183,
98'h071085ce0454d348a2d95645b,
98'h38fad331f05018a09a52baf49,
98'h38e388b1e49fe9093760dc6ec,
98'h211945020eb09bdd6bf27837e,
98'h235f5c86870a84ce0a9a78552,
98'h2b0168162a169a94354600aa9,
98'h1490f8e90cb0f7d948507c309,
98'h00dc0e41aa84e0152ad83b95b,
98'h39157c320919ce52308bd2a11,
98'h1f077cfe36a24cad756a726ae,
98'h106bb560d367b8e6e8f4db91f,
98'h160594ec3f77e0bef55f5d6ac,
98'h2613698c230e3106324866a49,
98'h28daba118c3883d86d44cf7a8,
98'h0abc5cd545e2e5cbe427d0a85,
98'h3bc77ab7ba748b34dd8f017b1,
98'h1d371a7a4b15de562a133e342,
98'h1876f970da8b04f50cc07f997,
98'h0fc97bdf9aca6775aaa4f8d55,
98'h306c1120d41abbe81121b3423,
98'h17f8f2efc8bab6d1682cea705,
98'h08a742d16ea5041d4dd311bba,
98'h18cc8ef18d80565b099339532,
98'h062f58cc73843fa70e6ce61cd,
98'h35f8c7abe1cb4b03b5f104abe,
98'h3656d02cbbc827b7bc87bdf91,
98'h155703ea8501fc4a0696400d2,
98'h134802669a79d474cb7075b6d,
98'h3f7adf3ef173dca2dc3baef86,
98'h39920a330e3984dc51f2e3c3d,
98'h0c2736d86f78d21eeee8023dd,
98'h32206f24781826303a8e25552,
98'h2fd4ed1f8a875cd52e97127d3,
98'h29378a125cfe9f79d18d8a630,
98'h106d7560eb7b8016eefa3d5df,
98'h12bfafe56ee4d29df06920a0d,
98'h1ccb17f9b5f86babd4b0e0e95,
98'h225918049f8a6cff3078e140f,
98'h3880fc3107fee04fd01ff7203,
98'h0e62865ccb5366d6866d7b4cd,
98'h3fdcf2bf8e825add3397d3673,
98'h1c4caef8bc5a5238b629c04c5,
98'h3304f8a613f6fb67d1befd037,
98'h1e44627c97ba5eef6d7fb05b0,
98'h168283ed2a822b1530412bc09,
98'h226d7504d583246b2dfc265c0,
98'h077d87cee6a8090d6b8964371,
98'h0698664d2ab828954c5423b89,
98'h3e593fbcb4ff8da9fcd63359a,
98'h3c8cc5b9282e2890792ebb926,
98'h3f54b63eb9a774337e3f0a9c8,
98'h36b261ad7d0820ba3ceea099e,
98'h22410b8486e5e3cdca49bbd49,
98'h3f13293e2406138818c64f318,
98'h244f80889d8cd57b10771580e,
98'h0f5fd6de83c79447a4c9dac99,
98'h3d693cbac16d3dc2cfb59e9f6,
98'h2bd157978f940b5f2ed958bdb,
98'h3172d522c252f4c4acf17279e,
98'h3070f5a0fc2ac0385b26ed764,
98'h294d97129ab35cf571003d020,
98'h3c813bb93e8ca33d1ec377bd8,
98'h03588fc6bc68cbb8cff056dfd,
98'h1e71a07cc5a1d1cb4904dc920,
98'h1ba351777d84b23b364a00eca,
98'h1ff6ecffcf0ce15e2bc0f3978,
98'h04f47dc9df7283fee919c0723,
98'h019266c3176de5eec640132c7,
98'h29360e924d555eda8da2db5b3,
98'h2301b48612c73a65ad723bbaf,
98'h05c95c4bb7ba752f4f60f45eb,
98'h2ec18a1d8ea6095d6f59e4dec,
98'h12b4e5654f6a335ec887c6310,
98'h2dfd0c1bf920933279c767d39,
98'h168dd86d1b522976ac780078f,
98'h1bf3fc77c1ac38c347680d4ec,
98'h106f59e0ea31b1144ea842bd4,
98'h30119ca03f3d413e5bd3b7779,
98'h39418eb2bbe35937fd4939faa,
98'h109e5d613612622c31ac2fe35,
98'h020261441bcd09778773daaee,
98'h01263ec25afe08f5e70911ee1,
98'h21b20c835230ede46cf8be99f,
98'h135dfe6685ef61cbc653580c9,
98'h16f560edf8c91cb1b3ef9f67e,
98'h3380fb2705ed1fcbce5b86bcb,
98'h336fcea6ec480018b7edf3afe,
98'h05d1e0cbb1a404a34ddd795bb,
98'h35472d2ab4077c283a53aa54b,
98'h3e180bbc3d1b2a3a3ecccd7d9,
98'h1a3342745760d8eeec6506d8d,
98'h0fa3b55f4b10085626acef6d6,
98'h12eb0be5e0d76881acf09d19e,
98'h1892d8f13aec3db5f4dfc5a9c,
98'h09b1c4d34e6ff1dce6086dac1,
98'h29c0dd139737196e503dfda07,
98'h2735b08e503ed3e06ddd211bb,
98'h11fafbe3dfd4df7fac73f6d8e,
98'h21e2a203c666f2ccea1265343,
98'h0ac36955b355d4a68f864f7f0,
98'h093a41d25a735df4c8eb67f1c,
98'h1b1d3d762f07039e328910451,
98'h24b418096125b58251767362e,
98'h258b1a0b3a66c734d7fc784ff,
98'h00175440158357eb0566ab0ac,
98'h2d9a961b340f1028386a6990d,
98'h1a3053f4401b43c00692e5ed1,
98'h1b0661f618176ef00cc774398,
98'h3a33ec346a2ec3147918abd23,
98'h28a92f915660d9eccfc2825f8,
98'h301271a01f96d4ff13ea51a7c,
98'h302b6020662d370c759625cb3,
98'h106c7f60e7f0508fce1733fc2,
98'h2c8563190fd4a4dfaf1681fe3,
98'h11cb7ee393c8d36789651492c,
98'h0920e6d2615a7e82aa9ed9554,
98'h2a2ff2146936619274d994e9b,
98'h2d92b99b2b1427161629b82c4,
98'h25f7788bf073d6a0f59ad3cb3,
98'h1a9776f5328391251346c2068,
98'h078c99cf08cc06d1a41628283,
98'h282ceb905ef7857dd1c91c438,
98'h0e424bdc944da968a8a3fd515,
98'h325240a4b973ac32daf17b35d,
98'h262d3b8c597200f2efe7cf1fd,
98'h0e28e25c4bd254d7a67ecdcd0,
98'h36bcd5ad411043420df3463bd,
98'h27e0260ff601fcac177888aef,
98'h26460c0c80a7c14149bb73537,
98'h3705b62e0fb099df51ad94035,
98'h31a1e2a3593ace7272b72c457,
98'h3684b7ad1ca69ff954cad5e99,
98'h0471b148c5a468cb628586851,
98'h0bcdb1579683c9ed08945ed12,
98'h0c8b30590c82a2d9064374cc8,
98'h31513622937fa1e6f13436026,
98'h2d7e3e9ad57fc8eaf0bf81e17,
98'h17a74bef7b3fc93654b9c5496,
98'h3c166b382bf44997fa02ad340,
98'h326d9324c4c600c9adcce4fba,
98'h212a3a026d8b611b33ad66c76,
98'h16162f6c3ee7ee3df53f876a8,
98'h2afa3015cec47cddae6fab3ce,
98'h16916f6d23b2a8876e9105fd2,
98'h08d198d18cdb64d9856b3f6ac,
98'h07ec344fca8bfd55049e0c693,
98'h298b0d1320d1240192970c452,
98'h05ad1b4b70d377218da0249b3,
98'h170abf6e3dffb2bbd5429c8a7,
98'h07ea63cfe1352a824a47e3948,
98'h2ab07e9563d2598793a0b6073,
98'h39c298b3bad039b5bd24b49a5,
98'h353382aa79ecdd33fbc817f79,
98'h0811f75016c31ceda7b5450f7,
98'h2b49f1169c3b65f871e155c3c,
98'h24ee9809c89fac512b639116c,
98'h33ee27a7d51524ea3240d3248,
98'h10a5576150b8e76168578fb0b,
98'h1103c26212cbc16588f3e0f1e,
98'h07a17b4f4a2c7c5464737de8f,
98'h238e640717b17aef4ecff7bd9,
98'h09d91d5385fa0fcbe3f4cb47e,
98'h3d9c3f3b03d01547b05b1520b,
98'h380852301c6a4678d51ca62a3,
98'h29765c12d23a7fe44eec36fdc,
98'h093511d262778b04eaeb2735d,
98'h0398a44705133b4a022af7e44,
98'h0ba5de575dda987b8a601db4b,
98'h1763a56eef11851e119d4aa33,
98'h0ba52dd763ccbe878bdc7b17b,
98'h196a1e72db7f3c76cd3a56ba6,
98'h041b90c80081eec121275fe25,
98'h39ac443372598b24bb0173d60,
98'h353a9aaa73cc7f27ba41c6748,
98'h1802cb70296e5092f05c4700c,
98'h10228a60764cb62cb19bd0234,
98'h016bae42c9004452229afca54,
98'h1f9cb17f35fe112bd566b0aab,
98'h01dab7c38eabe1dd6421a6684,
98'h21b49b8344e44c49c9a639f34,
98'h1f9fc87f37f70faff5e5b60bc,
98'h3029fa206d0a2a9a174d092e9,
98'h3f64e03ec325884650a29a214,
98'h0a6546d4fdf3fdbbf21651243,
98'h1635e76c6c9bff9930b479c16,
98'h1ec92f7d8d17efda0af847d5e,
98'h2df4329be54c0d8a94d010099,
98'h3eeabbbdc8de07d1b1f230e3e,
98'h3407d0281f52d4fe94d6a949a,
98'h066a38ccc019f5c001a10ba33,
98'h0e108b5c25246a8a6ccd3d79a,
98'h12d6dc659ae09775eb6ddcf6e,
98'h20c8b781a94e00129285ade50,
98'h08372fd0510b41e226509c6ca,
98'h0e3bb75c6508c88a2cd11ff9a,
98'h2d80389b2aaac915560ac06c1,
98'h0de2435bde87a2fd2b1a79964,
98'h3a755db4e31c48863764698ec,
98'h1f2673fe591980722e0ffd1c2,
98'h291b12121c61aaf8d15f2f42b,
98'h11418862acea8d99cf8b057f1,
98'h0c163bd809cfefd3a5798aeaf,
98'h2e556d9c9e5e1a7c932ce2064,
98'h3d025a3a131538661405e4a80,
98'h1f140afe31ab4123742fd3086,
98'h35f871abc7088bce0f403f5e7,
98'h143642687296502531b324a36,
98'h0430b14844a55fc9623584447,
98'h0774c04ee5d0ef8b8b516bf69,
98'h02d8d9c5a404e10809b76eb36,
98'h32a47e2565bb0a8b7617e22c3,
98'h20e96801dd16fd7a0f80195ef,
98'h0d090dda32ee78a5effde1a00,
98'h26f37c8dca4d2654ac5028b8a,
98'h30de9e218e2f635c4fc3805f7,
98'h2e91809d2e58de1c973a97ae6,
98'h198dc7f3310b6e2212a64d854,
98'h105492e0b18ffea310792460e,
98'h31eb1023f8a1a2317aa32c955,
98'h22b8ab055978bff2cf0c5abe0,
98'h0554344abebd10bd710451420,
98'h08d985d1a76f800ecc1241781,
98'h126d3064fc9c40b913c25c477,
98'h2e52491c8e484edcaf26a5fe5,
98'h16af076d546f51e8cac796558,
98'h32e1eea5e63e300c564807ac8,
98'h2aea4b95cec6e85d8e6c4cfcd,
98'h201e6b002e72281cf3a424c74,
98'h0e4f66dca3ddd187ac8b4e191,
98'h19b096735fac02ff6e57265cb,
98'h037e9fc6d9d771738755844e9,
98'h3942d23290fed961f2906ae52,
98'h0591e6cb04bce2494293b2451,
98'h3e7c753cd0635ce0f3b7f4877,
98'h1602596c1732e4ee4b4d4f969,
98'h1513efea1349de668a1773942,
98'h13bb8ce75f9283ff2cd38439a,
98'h3b31b536619614031731f24e5,
98'h2b9e9517103e7c606ef7445de,
98'h350de42a1466a568d25d2264b,
98'h1f26cdfe77bf672f55b98d4b6,
98'h03e2aec7cd7a6ddae4574728b,
98'h12d260e5a160a002ed0cc03a2,
98'h31fd80a3e7f58a0fd67cc2ace,
98'h2f608e9ee5b7ed8b75461f0a9,
98'h3fe8eabfebb81d975ae84215c,
98'h1ae7b875c7b1e9cf68a668915,
98'h035946c6bd68dabad03088605,
98'h053524ca426d28c4c1e89363c,
98'h23b622877ac54a35979edb2f3,
98'h31d889a3b25e2224b90daaf21,
98'h3dca66bba8b9d39159a10e933,
98'h2dad541b74e5d929d8a4cb514,
98'h24553f08ab33871653e23187b,
98'h31a3b12340b542416c963cd93,
98'h19e5c273e98da21330dcd921c,
98'h34fb5329c3076f462e00b09c0,
98'h0d9b59db21ecda03ebe20cf7c,
98'h1a11fc7405ec734be7ff9bf00,
98'h0414e9c83dca633bb077d340f,
98'h0e57c5dcb68f0cad1139b4a26,
98'h3408ba281660b86cf29a5ca54,
98'h23eb2787db8f0df70fde8d5fb,
98'h26af1e0d7c9c233918d2d0519,
98'h35cec12b973a82ee534251067,
98'h2b59db16a1a10603533eb8467,
98'h0a9ae0d53b9f9ab7318e9ee31,
98'h0f42515ea6e9e00ded8b0c5b2,
98'h00fccac1eb2151964b0787160,
98'h1ac86475836f18c6e78ddf4f2,
98'h1945c4728b68d3d6c92ba6125,
98'h000c23400a3a86544291aa651,
98'h03bbd7475e3daafc687e6090f,
98'h37fc2f2fd238b5e4728d39451,
98'h384e5eb0affea11fda133ff41,
98'h2ea2e51d4309f3462c6b3618e,
98'h1dc04bfba2256e846ff96ea00,
98'h21ac45037b0511b6372c55ae6,
98'h284a2e10b56f1caad76e52aed,
98'h20ce98819b8df3772f1722fe3,
98'h3625fd2c46f32f4dcf464b1e8,
98'h02efde45e651d10c8a506bd49,
98'h07669ecec1a38ec342428b648,
98'h0891ee5133eb43a7cf1f4c7e3,
98'h19ed3073fe5f2d3c9613176c1,
98'h183f64f046e009cde7c7dbaf9,
98'h2e3e0e1c7bf17037da8bdf950,
98'h30634720d0da91e1904f76409,
98'h22679a84ea085894131bfcc63,
98'h1f25707e4771404ec9a5ac334,
98'h211cc882025b6ac4a8de0cd1b,
98'h3895b4311dbd7a7b7594cbab2,
98'h389560b105ed53cbefa0ad1f4,
98'h299fca933c7469b8f9850d130,
98'h02b60bc5758256ab0e0e189c1,
98'h16f1f66ddf2389fe4d85601b0,
98'h3a721834f0156f203aa1e1d54,
98'h3e306cbc6ea2eb1d7b34d5f67,
98'h2549040a94463d688e63d05cc,
98'h397f7eb2c2bf3e456f0faf3e1,
98'h3731c52e7e69abbcdd66dc3ac,
98'h1d9e7ffb038d99c7084b06708,
98'h0735cf4e501757e005d349cb9,
98'h1d7d6e7ae9cb039391d21c839,
98'h276ddd0ec3bdba474acae5d58,
98'h37675c2ef919b9b23c2045784,
98'h3802793032f70ea5dabe61f57,
98'h1b8b96773ade3835959a73ab2,
98'h364244ac9508fbea32d2d025b,
98'h05df8b4b98ee0171c7b3632f5,
98'h12d00065a028fb004cbe3ed97,
98'h1a0376f4383227b0748d67a92,
98'h205a51808fcf81dfac0a74d81,
98'h3b03c63638cf94319cf4d699e,
98'h2b3f50166893e69114f4cda9d,
98'h0681424d07570fce83761486e,
98'h1dedc8fbd2bb0d654c2a35984,
98'h16f9f5edccef0859c8fa3f91e,
98'h39c646b39bd2ca779566444ac,
98'h279cd80f07591d4e8bbd7d576,
98'h3cadde3949640e52d1847b230,
98'h31423322812562c26c99e5794,
98'h0474b148eef5cd9dccda9fb9a,
98'h07d2cacf82556cc4828a0de50,
98'h3ea2383d5c4aa6f8b6bb37cd8,
98'h2d97c71b3e2117bc7aee37b5e,
98'h31294ba241f34b43ecc725b99,
98'h2a9d5a15377f0c2ed8871990f,
98'h02f5eac5c5ffa7cbe23d64a47,
98'h05822acb2f830c1f2d414dba9,
98'h1e36c3fc7cc8cbb9b6bfe3ed8,
98'h2cbd78196a93f81515d45c0b9,
98'h2db47b1b7e7d91bcdb0c83360,
98'h3f9606bf0feb965fd3e06747b,
98'h0e78b5dced4c071aaef12f3de,
98'h20b3c50155c21d6bad9d789b4,
98'h3376dea6ddb195fb744a1d289,
98'h1d6634faeff77a1ff3576bc6b,
98'h25d8af8bbeabe83d792125f24,
98'h28699290cafc58d5ecd97ad9b,
98'h1e007a7c063494cc690d43d22,
98'h3924bdb25d2cecfa55946aab2,
98'h23432e0693a186676db92d1b8,
98'h3d09e0ba01bf77c36fb2561f6,
98'h0ecc22dd993420724a0010d3f,
98'h3bf3da37fdd893bbbe731b7ce,
98'h350c9daa3c512b389c577238a,
98'h060a61cc3e4737bc911466622,
98'h34891ca9248b79093645256c9,
98'h05e6f34be6da830dab305d966,
98'h34c65ba9b0db4fa1b9686ad2d,
98'h10647560ef33441e6fe5ee5fd,
98'h18881e712c0c8f9811252b824,
98'h10b3a1e160634080ec45b8989,
98'h0783b54f299d9d130c4854988,
98'h26fe2d0dce9c3bdd2d669a3ac,
98'h19184b721ef905fdee04545c0,
98'h0612af4c3ea0c13d712cdc226,
98'h0f8ee75f1e23ec7c6b6cb4f6e,
98'h3d434a3a8398aac71036fd406,
98'h15d4396bbaab2c35541fd9683,
98'h32d11425a35b6986958b1f6b0,
98'h0c8e1ed923c945878c15d9182,
98'h0cee3dd9f1320da26f8812df1,
98'h02deed458b6f03d6e3937c472,
98'h2f90fa1f2d830e9b3745022e9,
98'h371878ae1508e36a130857060,
98'h380128300fc9d2dfb1f2bec3f,
98'h0810dc502c8b3d190d27065a4,
98'h083ab9d04babf65764f9ac09f,
98'h14bb02695a7f2d74ebce8bf79,
98'h2feedb1fddee55fbf3774c46f,
98'h0114eb42187a3a70c663c96cb,
98'h1b1ddbf6167bd46cec666c18c,
98'h316db7a2de9abd7d14021d47f,
98'h12f3d6e5e59fe40b0e24eebc3,
98'h23756f06ca530ad48b721e76d,
98'h18c219f18806ced008323a306,
98'h1b788776e4fd5b09f01d78a03,
98'h209f4d010305bb4628e94211d,
98'h3f992cbf21627102f83ee7708,
98'h3d685c3ad51c79ea34a135894,
98'h2ec84c9dae8d019d1755538ea,
98'h168c1e6d099307d32807c9901,
98'h01b059c367f3dd0fea690db4d,
98'h0d3bbcda5d84dafb0ab025f55,
98'h2cb3d5994334d8466bfa2b77f,
98'h3649dbac949be6e912b970a56,
98'h07919a4f0e4a715c857702eae,
98'h0c3283d8582d66f04917fab22,
98'h0d30df5a6a5638948de1c5fbb,
98'h2575c60ac05a654089740ad2d,
98'h108703e11ac9fcf58ad44035a,
98'h1a9f2a75104602e0aab94b557,
98'h2679160ccae9ac55ec58b098b,
98'h0903cf5238637fb0d059d3c0b,
98'h3c0b1bb8005001c08f16c75e2,
98'h0f7159def84e03b0b1efd763e,
98'h381f17b01c4feaf8b51bc0aa3,
98'h2cb79719788c24311950eed29,
98'h3c75d638fbbcb0b75e0ca1bc0,
98'h1926eaf248112e50284e0650a,
98'h169370ed00d2dec1a5d993ebb,
98'h37cd6faf8d3e2eda5142e7a27,
98'h1299986509abeb53471160ee1,
98'h1e6ce67cca94b8550a4067b47,
98'h24199d8812d69fe58dbc0f5b6,
98'h1fd3597f903d6ce06c0431980,
98'h175037eeb55e41aa932b9e664,
98'h077085cef0f445a1ee1932dc3,
98'h342d0ca85dba77fb7479e128f,
98'h3ab204b54edc9b5d9263a804b,
98'h07f7f94ff1d1f523ae727b9ce,
98'h08e031d1ef2eec1e6e03c77c1,
98'h2656198cab69df16f46ffe28e,
98'h00e5d341f6a2672d4de20e9bc,
98'h3ae09135de0bf77c163b222c7,
98'h399c833317e430eff4602d08c,
98'h356f122aff9d7fbf1d43247a7,
98'h00e7d641d55e6dea8591910b1,
98'h10a825e14590e84b058e438b1,
98'h2c1943981c010878320693041,
98'h2859331089cc31d3ac8959391,
98'h34c6cea9a9ae3b93579d428f3,
98'h27884a8f1e0e197c11659902c,
98'h346e6ba8c35cd7c6adf2d0dbe,
98'h0121a9c246cbfe4da1fb6a040,
98'h1af02cf5f0f24da1f2f89ea5f,
98'h059305cb33328ba66e31645c6,
98'h341924a82346740695d7e62ba,
98'h379692af3b231eb67cae6c596,
98'h232912064fb3115f6cb708d97,
98'h1edfcbfda1b7f0035025ef003,
98'h346cc728c80122d02f1b7a7e4,
98'h3c4bfab89f08fbfe16d53dada,
98'h30b750216175e382d48b4ce90,
98'h0ca881d9729ba8252fd10a7fa,
98'h08b3dc51763197ac6fb95cff7,
98'h3110dfa205172eca0d8a039b0,
98'h22ba67056d02111a33ef1e07e,
98'h3a567c349787c46f34779028f,
98'h21011d02193af8f24e8f057d1,
98'h33d42da7b4aa80295a1fab743,
98'h03b488476a15d7140b7297d6d,
98'h3d7f813af96c0532fdbae19b7,
98'h26b0728d638bdb07328f13652,
98'h08f9c2d1e0f3e901ca7b6af4e,
98'h31439422b58b62ab19b3bdb36,
98'h3dd2c53bba46dcb4be06687c1,
98'h2b97f61715db436b905cce60a,
98'h221f6a8415b992eb4df63f5bd,
98'h3d0a1cba00edd0c1cf7dfb5ef,
98'h01f5ecc3fb1e6b360f4515fe7,
98'h24e8f009d255a6648dcfa59b9,
98'h2e51e31ca2c7d605b4466e489,
98'h37c862afba7e2db4dc91a4191,
98'h26520d0ca729818e535ee3a6b,
98'h1ac0d9f590b9e9616adeb0d5c,
98'h10b1d9617f123cbe13f10587d,
98'h07a5564f5aa877f5689373913,
98'h32d0aba5b528a1aa79fe53540,
98'h256a5c0af86660b0d7742f2ee,
98'h0a88e9d50c847ed905c35a2b8,
98'h1aa7997573e89aa7f3a40d075,
98'h3488bd293feefbbffd1dee3a4,
98'h014e50429555d2ea85a908cb4,
98'h15cea16b9583856b2ad489b5b,
98'h365e7cac921f74e4121f7c642,
98'h305ba6a0871b714e0dddc5fba,
98'h3294bea50d0c735a0fe84c7fc,
98'h1d1d7dfa0d1e695a0a8ef9d50,
98'h15bb016b6657d18c8f04b4bdf,
98'h33823d27190192f21320f4064,
98'h2175e102e874e810d27ab244e,
98'h2e17eb1c0aef7455ee41d7dc8,
98'h3618d7ac2bfb6f17d88511b0f,
98'h3709c52e16c2a16d937319a6e,
98'h083b205077ad45af4ffa197fe,
98'h333d47a66bad1e9777ba998f7,
98'h24776108e477fa08d23bd6c46,
98'h3b40f4b6b3968e271bb5e0b76,
98'h3bf014b7c4c41149b02d09806,
98'h322edf246f6b121ef8667c50d,
98'h0be2af57f6540f2c908dafa11,
98'h3014efa00044fa408c167a782,
98'h08c38851ba653fb4d0ca32019,
98'h3b64ef36de8b277d367c05ad0,
98'h360c82ac2cb43c1978b02fb16,
98'h2f5e4b9e83ce3647accb20799,
98'h0b1873d613773666e7a3ea8f4,
98'h2853a490ae5e669c95ac82cb4,
98'h1f154bfe044ffdc8a8d95271b,
98'h3e1e0e3c124443e4941894882,
98'h1e46ff7c98a7c9f16dbbb25b8,
98'h35001c2a0e760a5cd0dd89a1b,
98'h2d852c1b22d6c0059416fb082,
98'h39aaab3342d3d345af1f9f9e4,
98'h2a0d849420e93e81d2bdb0c57,
98'h320563a437a47a2f5a6a7774d,
98'h0f74f55ec5c4e14b854e75aa9,
98'h05cd07cb95fd466be6f2938de,
98'h07b18d4f79df4b33b0643620c,
98'h3c0977b805ae504b506df200d,
98'h2de7271be5a8ae0b74e3f549d,
98'h00cd79c18cfdad59c372c9c6d,
98'h27d0d08f8d3c135a4d4338fa7,
98'h15a244eb54ab54e94a9366752,
98'h1750f36ebad76335948a15a90,
98'h3270c5a4e367c906d57623aae,
98'h11e239e3c80d2c50267bd98d0,
98'h30aaa8214b1780d60ef08a3dd,
98'h32533a2480922d410cb959d96,
98'h1ae52075cbed0bd7c9b48b136,
98'h0666dfccf8f89b31efd7debfb,
98'h24076f082993fd933366db26d,
98'h39a38db3439b2a470f4fadfe9,
98'h369f2f2d015695428dfd711be,
98'h3ccb0cb98a69d554d1cd38839,
98'h3adc5735a9582412b90d1ed21,
98'h32252ea4793a66b27ad7e555b,
98'h3c2706b86cae36997a354f547,
98'h25f7390bedaebf1b74e97e09d,
98'h3a310bb462527d04b720e22e4,
98'h3c320d384bb2df5751f93b23e,
98'h08d52c51919771e3069b278d2,
98'h0c910ed93c04ae3812256f444,
98'h2a062b1421f9c203f2fffb460,
98'h1113cb62392781b2728ed3452,
98'h217f9482e1d87683b0d602c1a,
98'h1bec65f7c295674507a0734f3,
98'h1eda427d8bcddbd7aaaa07955,
98'h2dacb99b51f02a63cfe738ffc,
98'h1c16a57809132752294a73329,
98'h06ac474d5e641efce94419929,
98'h309ecd210c88e2d90f49ebfe8,
98'h1b50d976935ea666ababdff75,
98'h3732322e71ae13a35a3811746,
98'h3613ecac3d2a7a3a7ccf99b9a,
98'h3c1d3a38190020f2354756ca9,
98'h37cedaaf8bf3b2d7f0f0a361e,
98'h148e81e933ed7d27d21effc43,
98'h1b07bef608258f5048cb53919,
98'h3bcbe537a1b50e8377603ceec,
98'h0da91fdb6603fc8c2ceb4719e,
98'h3b7947b6d03c556052ed6745c,
98'h29be56936dd2e19bb5e44e0bc,
98'h35131baa141654e8324a5c249,
98'h3d7eb83ae5cd210bb8d2f651a,
98'h382eaa3045a53c4b4f74f99ee,
98'h39217cb26f9d671f1a2fb8f45,
98'h27021a8e3270cca4d65cb9ccb,
98'h29a4669357faad6ff067c500d,
98'h1d263d7a457b834ae8a870315,
98'h2edf2b1d887a84d0cdd66bfb9,
98'h17740f6efb907fb734c123c98,
98'h04ed9ac9dd9b1d7b08a22e113,
98'h1b500676b5342baa54210c883,
98'h112a89e271770ea2f0a866215,
98'h0ba516574b11a5d625adaf0b6,
98'h15a576eb7284df25120a95841,
98'h16417a6c9f6ee67eed6c183ae,
98'h072cf24e79344b3250184f602,
98'h29373c924b61a8d6ed26395a5,
98'h2db7ca1b7b2b4f367a38c6547,
98'h09527e52a52f140a6ba064974,
98'h0126edc25354ee66851ef70a3,
98'h2ca77f19427021c4ebc5e8379,
98'h090a175216e3baede7fb74900,
98'h02aa67457044c6208cbbcb597,
98'h31413422b4da1da9b986d4731,
98'h1232cbe4720fd9241110a9421,
98'h33048e26239a5e8715a7bb2b4,
98'h293cf99257e5bd6ff048adc09,
98'h2e0db01c02706dc4cc1f87783,
98'h3e2afe3c7507c82a3cccb199a,
98'h044b10c88ff7685fe5109e4a2,
98'h32b76ba558766af0f2cb75a59,
98'h07b8794f45ace3cb43595746a,
98'h21bbe40371d41823b4e3ff09c,
98'h39a62f3348f3f451f0a688e15,
98'h1e5d617caf82ef1f33781426f,
98'h08e8d951ce39f4dc45c8b38b8,
98'h09203ad26c1721980d4dd71a9,
98'h151c2aea3fdf0fbfb53eceaa7,
98'h39d5efb39ce81bf9f5af82eb6,
98'h0c5248d893f485e7e811b3b02,
98'h3046aea0adba6d9b7780470f0,
98'h2a39f49475d2b72b98032aeff,
98'h24e89c09fa2c71b477c5436f9,
98'h3ff5713fdef8ebfdd7bb974f6,
98'h2ae6dd15f0bfb5a176e9a4add,
98'h268c2d8d2998d893340941881,
98'h392a5bb2490921d2308cdf612,
98'h1f112b7e2a9feb15126c45a4c,
98'h1d06537a22c1e205aff20d5ff,
98'h174826eeb500502a33121dc63,
98'h2a9a93150a230d546d2f681a6,
98'h1bc37ff7a86bba10d10bce821,
98'h30ed8d21cb260cd64f04e67e0,
98'h1d24e17a56a1eb6d4cf1b339e,
98'h2630178c5cf3c4f9d0c8f7218,
98'h215aa802b7e4fcaff64fe92ca,
98'h278cf88f0cfc7d59ed225d7a4,
98'h2f640d9ed51566ea111e5d223,
98'h23562e0699e28973ef4e2ddea,
98'h08560d509867c870e82f75706,
98'h1051f360ad91ae1b0f78e85ee,
98'h3f0b0dbe18966ff115e85f6bc,
98'h0d598b5a878d4c4f2539b5ea7,
98'h0517484a09e0a1d3e3bdfa878,
98'h256bc88af8af47315786c3ef0,
98'h3b4bf1b68819a35030d96541b,
98'h19c55473bc41ae38b581c0ab1,
98'h0a4321d481797e42c2ef2805d,
98'h3980b6b30b8d2257314376429,
98'h281e7a9026d18d8db3bc02077,
98'h10b01ee16ca600196f5587beb,
98'h07d292cf8736c2ce43c255677,
98'h13d2ea67bf72483ef4d14ca9a,
98'h28091a101f23ad7e51cb31e39,
98'h3bf8eeb7d89243f13522ccaa4,
98'h1fd3c47f8184444308560230a,
98'h07d5804f9d05f17a2936dc727,
98'h0a19f0d4180d6df02889d7b11,
98'h22743984f719292e366358acc,
98'h19db0ff3a3b247074f6355beb,
98'h0531854a715087a2ada0833b4,
98'h1d0fcf7a21f92d03cfc23f1f7,
98'h2408e48832c1122595b27dab6,
98'h0e23fe5c64628188eca19ff95,
98'h0d3af75a4d6ca35ac6a9e6ad4,
98'h38b33731780337b01c2d9bb85,
98'h3bbd443776ed0f2ddcaa94d94,
98'h31624822d0e517e1d091d8012,
98'h2ad5c215a9e80d93f52f73ea6,
98'h1e5f597c82aecac5684389108,
98'h1cb41e797f75e13ef70a7fee1,
98'h1a42d6f482859f4507321d8e6,
98'h39cac43396d4bfedb427e1085,
98'h01bb16c3790b13322eb18a7d6,
98'h0f19a6de0b72f9d6e6a3282d4,
98'h099cc2d32ac81c15ad1937ba3,
98'h3a8cc9351189e2e31305ab060,
98'h3aa200356d482e1ab9fa8b940,
98'h2200838404337948698cff332,
98'h2e52559c9b960477127a1684e,
98'h1f6d8efec914cf520a2097943,
98'h113d56e241bc284344be5fc96,
98'h372ec92e59673172d4257ea84,
98'h0de2085be05b3b808b8f50f71,
98'h3042c1a08a5a0e54aea733fd5,
98'h054d0bcab357ff268e2942bc4,
98'h1ddafcfb8377a1c6e854a7b0a,
98'h2aa783956d13189a35eea70be,
98'h117afee2fce65939f39856073,
98'h21a0bf83568c9f6d2e0b57bc2,
98'h215913028d10fd5a2b9a84173,
98'h30cca0a198455ff0924480248,
98'h2ba2d397496f98d2ed449b1a9,
98'h1cc0c3f9939fe5e72c182a783,
98'h20b7718174db23299564a52ab,
98'h22ea6805c4f34549e9f76b53f,
98'h2059bd00b305e62634d7e8c9b,
98'h37c7192f9f71a07ef5ce2e6ba,
98'h344bed28a862a590f72ba4ae6,
98'h2f5a139e91746f62f033a0c06,
98'h29b727935bf48a77d16aec82c,
98'h3c6870b8ddb08afb76863eed1,
98'h1630ca6c4931c55247d8a3efa,
98'h07360bce5043f1e085de7f6bb,
98'h311f70a21f52fdfeb41c9ba83,
98'h2b2d2b96497f52d2ed2b1f9a5,
98'h32b1bea55d19737a33f2cc87e,
98'h000ae9c03fbd523f6ff20effe,
98'h1a88e5f51845e9f08cb3b3f96,
98'h1ada5af5b18994a33318fbe63,
98'h35a8eeab7aaa50357c14cfb83,
98'h3938763265c9858b97c07eef7,
98'h3130c2a25ff027ffd4483aa88,
98'h3a0abeb40488dec92fa4e75f5,
98'h19cbeff3b2ddada5932a67664,
98'h2e02aa1c247bf108d49fa6c93,
98'h12c034e5bb13c0b63374fd66f,
98'h13f7c967db39ad766bcc5db79,
98'h2ee8c69de8ee8b91d5f5d48be,
98'h0d52af5a8c9f69d9267c864cf,
98'h25e1598be062ed00d19111a32,
98'h29729a92dcc06cf9918cc1e31,
98'h3c12e8b839629cb2fd5d615ac,
98'h2027dd806333338670d6c441b,
98'h19443e72b081162112715524e,
98'h1f0d047e0a7e7ad4ca62dfd4b,
98'h12c03ae581434042a500deca1,
98'h37b8beaf7ed8053d9da430fb3,
98'h1813def028b3d4917031ece06,
98'h31728722f057242098726ad0d,
98'h17d611ef8686884d2797268f3,
98'h0c440bd8922d0264479c438f3,
98'h10db29618943f252a687c6ed1,
98'h10f15461e664a60ccdd57e9ba,
98'h37a632af72a835255a9399f52,
98'h2591ad0b281cc010136b9b46c,
98'h1bd9f9f7988e67712d1a185a3,
98'h35334caa411d2dc20d941e9b1,
98'h29dbd2138072b8c0ca93a2b51,
98'h1623bc6c471a444e074f802e9,
98'h3dca1dbb9bc55d77b663deccd,
98'h2a2701147ce7d7b9f9c3b6339,
98'h1a5895f4adf8331bf21432442,
98'h02178244204e0300a89961513,
98'h341452280e612cdcd09d5fc13,
98'h0718b2ce2221b1044a4e98f49,
98'h3c0192b833bb76277bef4237e,
98'h1ab678755fb2e27f4e9a56bd2,
98'h2775440ed1415ee28e2da8bc5,
98'h30fb52a1ce92b6dd2fe3825fc,
98'h3a7c4d34f20901a41b2153b63,
98'h27b7460f6223360452769f04e,
98'h121290e43a7dacb4f3240f664,
98'h38e181b1c152d6428e8d15fd1,
98'h2fdbba9fb580082b3956f0b2b,
98'h272ec60e4655c3cc8b612276b,
98'h15ffc4ebdee6ff7dcd39b11a6,
98'h17a690ef761eebac33715f26e,
98'h333d402663cb690795c22a4b7,
98'h3d31013a7dcac0bb9ebef07d7,
98'h31335ca25e386ffc73daf327b,
98'h37c7812f8d1dc4da313951827,
98'h0555b24a918ab6e325b81a4b7,
98'h1c222f7872a8d12573b2c0277,
98'h2bebc697eaf84695f5b9034b7,
98'h2e6c039cec151e1816a0486d3,
98'h0fee56dff26b3124d09662012,
98'h3eb7ba3d478a0acf119071431,
98'h0e845edd3708fd2e31635702d,
98'h349f79a9360ea52c3aab87b55,
98'h1d51e1fa8470ca48e870ab10e,
98'h3ca93b396638f28c78b88b717,
98'h1bba72775dea3cfbee692bdcd,
98'h21b9f383666cf68cf209ba841,
98'h1ca97979476f224ec90626f20,
98'h33117aa6025d7d44ad5bbdfab,
98'h3c623e38d5a9ddeb548307090,
98'h17f932efcc709fd8c91a74b22,
98'h3849b13081b28ac34e7f0efcf,
98'h297f7192e51a0f0a13a660273,
98'h398befb31f84e97f3644364c9,
98'h0449a848942d1ce8661db14c4,
98'h32ef8f25c2d90445ad7224dae,
98'h0cb749d946987ecd04d3f2299,
98'h1218a3e4213898826cd44f19a,
98'h023f74c479eddbb3ef0b541e1,
98'h30ed8821c5db3fcb8db231fb5,
98'h08235b506a8710150caa9ad95,
98'h28bf6711400354c00a30aef45,
98'h253f690a750b38aa1692a86d1,
98'h0248814483459e46a16387e2d,
98'h36f52f2de485780916dea9cdb,
98'h378236af0655b64c8f75fb3ee,
98'h17d8076f972f816e4bc1e2377,
98'h32c4cf25b4a1312979d98013c,
98'h15f67f6bd981dcf32bde1717c,
98'h2593000b0d3386da6cb1a1b96,
98'h324a7f248d0bf25a2fd59c5fb,
98'h14e336e9fa0cb9b413bbfc277,
98'h0f0a33de0305d1c6248401691,
98'h0ca89fd95244bee4a7bb57af8,
98'h1943b2f29d7db8facdb05afb5,
98'h2ccded998305a7c62bf4e557f,
98'h275d660ea9735c92d43430a85,
98'h2ac3e295939687e72f969a9f3,
98'h25c5320bb422f1a8567a08ecf,
98'h103598604b611d56e6e5ad6dd,
98'h09485ed2ba31f2b470de9461c,
98'h2d64861afa0c3a3419dc3013b,
98'h073e3ece745fa9a8aee77a1dc,
98'h001e4bc02d74eb1aeb64cdb6c,
98'h12df97e58ecb78dda86ac430d,
98'h332e37264b805f570faba59f5,
98'h00d4c9c181d2dec3a0a9ea215,
98'h319c8d233a709234db0347d5f,
98'h0234b8c469f94313eb0b7ef61,
98'h10fd92e1cd95b05b27a4d0cf4,
98'h12de73e59b3b7cf66b867c370,
98'h2a82519539e64333f91a25324,
98'h08479bd09fa1187f69fa2d140,
98'h176d256ef23815a472694ec4d,
98'h11898de314cd61e9a995bbf33,
98'h06fbfe4de183df030a1ff7543,
98'h3ba749b74cc22c59b21a5d844,
98'h05ca6ccb96cda96da726058e5,
98'h19b619736ef6599df22b1cc45,
98'h2d1d679a05fbf7cbecc657d98,
98'h13c2fae7b45223a8920547a40,
98'h077ad54ecf17b35e25a4a22b4,
98'h04fec6c9f693222d2ee47a3dc,
98'h235ed286b61ecdac365f680cb,
98'h05eb194bc60a144c22fd4b660,
98'h08d0bcd1a4c3ac89ab651a56d,
98'h2df1f79bcb9468570e6197fcb,
98'h2f09f51e21235102540b51881,
98'h0d023cda042382c864496fe8a,
98'h20506f00a4ac3f09713f2b828,
98'h057abccadb13c8f60823a1703,
98'h0f96f35f192024726a2dc5f46,
98'h14de2f69ad05641a3078e4e0f,
98'h39652a32c2ca4345af0bdb5e2,
98'h2a79d694c9d8d0538d14a9ba1,
98'h1bf962f7f2b497a573ab7ea75,
98'h3258e924bde11dbbdc0e81b81,
98'h1d861afb0dd5c1db8ad6f735a,
98'h248eb7093c4dfcb8b8372cf07,
98'h36dd47adb2e1ac25fa6fbcf4e,
98'h01119442133f84666514462a2,
98'h28cb5d919b96f477311894823,
98'h13107ee618e5ba71cafd8e55f,
98'h3ed417bdac1312981ab9ca956,
98'h2fdd889f9c7ddc78f316d9462,
98'h26f2ff8dc6e7434dcb7690b6e,
98'h1136fee251ef66e3e8c999719,
98'h0f71b75edb582c768ab278f55,
98'h34e94fa9c73adbce6f090ade1,
98'h05d5fecb886247d0c38e11a71,
98'h0073b740f3dc4e27ad14015a2,
98'h18597c7086cd0a4d87c9a1af8,
98'h1289a2e537b3a6af728f52652,
98'h3a4d46b4a2c6cb05b745046e9,
98'h19fadaf3e4f4ae09cfbbe23f6,
98'h3f3b2b3e4e336ddc535ba646a,
98'h05bc6a4b5310d2e606334f4c5,
98'h2486b5090c07c6d80c239ef84,
98'h187c48f0f37cb3a6d2fe3f25e,
98'h31bff8a34ebbc6dd501eefe02,
98'h2759bf8e90a365616dff493c0,
98'h30ca17a1ac0d62181735de6e6,
98'h3b0c93363f497b3e9e95839d2,
98'h3c678ab8eafe3715d9d97073a,
98'h38f4ebb1f711d22e3c01af780,
98'h21ae2a037a25f7b456f5086de,
98'h123dfae47bc612b793810366f,
98'h2b54f516b823903078de2151c,
98'h066d674cda74fef4c83899906,
98'h20bd9a017227102474b92a897,
98'h386970b0f76876aefbf479d7f,
98'h2a0bbd94013e52426ad283f5a,
98'h352fdb2a60654080f56546ead,
98'h228c04050a3e63d46b3299f66,
98'h062795cc459693cb02ef8a65d,
98'h071cd94e01d3ae43823c21e46,
98'h0a2721547ef75cbdd2479f848,
98'h1b3af6764272dcc4e76b74ced,
98'h03f9bb47d7fb476fe6fd40adf,
98'h30c3aca1a894851136560c6cb,
98'h1f5d427e9ba987776ec1b27d8,
98'h306eeca0d6d592edb1d11fe3a,
98'h0a22e154444b5e48839b8fe73,
98'h2f730d1ee3466886b4ae5d696,
98'h324c76a49f40667eb4633748d,
98'h05b4544b4d62cfdac4c5c9098,
98'h2fb0ba1f637a9606d4cad4098,
98'h13523f66a4dc99898e0bb63c0,
98'h23e02787c3940dc709dd0d53b,
98'h30548a2088930c512e39e59c7,
98'h19b4a5f367609a8ef04550209,
98'h39a9f8b346c1084db01ac0404,
98'h3325ee26504d0360b0dcbc61c,
98'h0f9adbdf379bf1af11cdb3638,
98'h2bacb59773ce0a2797deafefb,
98'h3f415dbe964d566c9563ad0ac,
98'h2bae93976b913b9735cff3cba,
98'h368985ad2d61589ad8fab791f,
98'h0a1caad438117130308b87011,
98'h24ab03894f73d4deed07b61a1,
98'h309f10a113a11c6771100b422,
98'h03feb547d7164a6e26c53fed8,
98'h1056f660b5ec4c2bd190d0a31,
98'h1981eff33598842b33c69d079,
98'h3d718ebac664794cd0f58201e,
98'h3649872cbb8dffb73c75e1b8f,
98'h0a75b8d4d2f80965e75b708eb,
98'h139696e72b9a15972fcc2b1f9,
98'h2566660acbe798d7ec537fb8b,
98'h372f08ae5c3ce1f874dafaa9b,
98'h3483c3a9017b0442cd7fb1faf,
98'h070bddce1c0aeaf828c5b2319,
98'h0aa5205548c82ed1a4db53c9c,
98'h0d5f365a80e989c1c39230071,
98'h2fd5971fbdad8abb7b60c876c,
98'h046419c8f29a13250dbf8b3b7,
98'h360d762c2d92611b18e7f5d1c,
98'h1059fde0a70dbf8e2dd9ef5bb,
98'h0f9265df0c6ed9d8e7004fee0,
98'h317e0f22d7ac51ef524a98448,
98'h28b85091480dc4502c3185386,
98'h2bc43b17bde77e3bda6aee54d,
98'h0d6d0edad86a1e70c975cb52e,
98'h0281f4450f2515de4469c288d,
98'h3028c9206b7a5d16d6e8c98dc,
98'h2f2cbc1e4839ecd04dd9aa3ba,
98'h278d240f3aab7535788e26512,
98'h07be6ccf4b5f81d684c77ba97,
98'h362d282c54bda16952bab2656,
98'h17413deeacbe651950ffe8c1f,
98'h18a7e6f16ba4eb97511334a22,
98'h15758e6af557652a92b33ce55,
98'h356fe6aadf7f757ef53bd70a7,
98'h2d736c9aee45709cb6ee374de,
98'h0b4947d689a37e53653b318a8,
98'h3a99de351b0242761567082ac,
98'h2bb8ae1751372e624f3bf71e6,
98'h0b0de6563487c7290fe56b5fc,
98'h194ce7f291b41ae34ac040b57,
98'h2b7b5096e4d84909b414e6682,
98'h12dd5765af28909e70817a010,
98'h3cb937397ea7533d7ed8229db,
98'h1887187117f89d6fcc1fed783,
98'h35644aaae38d5b87163c698c7,
98'h1962eaf2c450d2c8876cef6ed,
98'h3370dc26c8602c50cef4421de,
98'h259dd98b3c6cd338f882ab310,
98'h0026a24076fa0a2dedc82b1b9,
98'h03cea247ac439818ac048e981,
98'h1fe8437fdae99c75eeb477fd7,
98'h0e11dd5c091b79d225cb55cb9,
98'h12989be53f3495be54734c68d,
98'h0fa6e65f67f7f68fcde7b73bc,
98'h055fc84ab2871ba52df9b8fbf,
98'h2a778394d6c33dedb04eb060a,
98'h3f01ebbe38d9efb1bdf6f6dbf,
98'h21244f827185732334aa70a96,
98'h00e9b8c1d1c95463a4acc3496,
98'h29dfde9384ebbc49ebb2e6b76,
98'h0c78b858d586b8eb087fdc50f,
98'h3492a82933d102a7ba18eab43,
98'h321f51a40b7f1e56cf679bfeb,
98'h3f71af3ec26a8244d0770c60e,
98'h222e9504518041e30cebb5b9d,
98'h3c61e838fb2a0a365de2fc9bc,
98'h2245c004bc5682b897a710af4,
98'h1332656653580c66a9a29c734,
98'h29ad8813778d8c2f384ec510a,
98'h04e73949e3d75e878a2fa5f45,
98'h36e3212ddd2dbb7a7504372a1,
98'h06ff22cdf174c7a2ee1cfa9c3,
98'h0d05065a340048a8304153c09,
98'h26cdf38dbb94453718988e312,
98'h2cc381198714304e2cf5ec59f,
98'h10b5b8e153fe1267e92cf2d25,
98'h25e6f40bc7edd8cfcb753336e,
98'h0138a0c27afd7235cf0d84be0,
98'h086dde50f1fb7b23ee9a565d3,
98'h1a8da7f51bf337f7cda037fb3,
98'h22b4a6855d984cfb10133ce01,
98'h2491f9892bee0b17f42001284,
98'h190924722718648e300862401,
98'h0aa120d551ca75e3871ae5ae3,
98'h167be3ecef07659e1160d262b,
98'h070de74e01cca5c38236a3446,
98'h1ab131754ff3e5dfcaa945d54,
98'h02a604c55195f963250eff8a2,
98'h18e3dff1dfd1957fae2d5d5c6,
98'h0bda82d798c845f18928b2324,
98'h353bd12a7b2c27365c19fe182,
98'h18d6e571b298df2512dbf125a,
98'h0b0a3f561b14fbf62987ced31,
98'h160114ec010560c205c19d6b8,
98'h046dc1c8dfe582ffe914d1323,
98'h3b0c0336274c340e98960dd12,
98'h065017ccb6a06a2d6f3c207e8,
98'h0ff7165feabadb954eac7c7d4,
98'h069fafcd18eb8171c7e2cc4fb,
98'h1d044efa02d3f645a7f6114ff,
98'h2a16ee140c4c62588d98d41b2,
98'h00df30c1b83f0b306e478efc8,
98'h3ed3383d8081db412fd544dfb,
98'h02de69c580e41141e0f09ec1e,
98'h2d6db79aea84141515fc72ebf,
98'h387a3cb0eb04b51638dfbc71c,
98'h0737e7ce45e579cbc34758668,
98'h28c1a5119d15637a3175c222f,
98'h09add9536cfe6199edab0ebb5,
98'h0ac8435590880de106d4144da,
98'h01203c42457d75cac1a76c834,
98'h38b701b176aab82d7bd86e77b,
98'h030827c63ea6db3d506bc0c0d,
98'h04597dc8842bbac842214e243,
98'h3f66a1bedcbc18f97708aeae1,
98'h2fb2301f6dc5cd9bb75dff6ec,
98'h0401e7c835b6c1ab6e6e2a5ce,
98'h304f54a08b05d0562ed5493db,
98'h38427630a2afdb0576bc944d8,
98'h02ca91c5970c50ee0675b8ace,
98'h30e1cf21eafe0695d6f7f56de,
98'h390d61323e9cd3bd1dea8d3bc,
98'h3b8d05b71e4466fcb6745b2cf,
98'h05a437cb52bcdde56618456c3,
98'h080d02501d5c4afa895a5352a,
98'h1c9a6cf92b94ba17120bc9c40,
98'h1a768df4c33393c6476a886ec,
98'h0308e346043402c841cf39839,
98'h14541668a269de84edaf7d3b6,
98'h1db1707b794be8b295bf564b7,
98'h1dab3b7b6ea66b1d731469a63,
98'h28b1041156e13c6defe4901fd,
98'h2630108c5550c46a8ee0353db,
98'h0a8293d51f68347eea7ab2150,
98'h16e82aedcc8626d928db9471c,
98'h173cbcee6dabf69b513a2ce26,
98'h38ef65b1e4d5ab89b771444ee,
98'h222431045e53e17cb01e04a04,
98'h0b006a563e7d2ebcd25f6644b,
98'h175cddee89c88fd388495b708,
98'h18d2fa719190f6e32a98fc553,
98'h11b3d1e35faaa5ff6c579df8b,
98'h2151f6028da81cdb6bbe84b78,
98'h252be78a65fd548bf2ca4f059,
98'h0f1b245e1d57b5fa8b1cb6962,
98'h32272d245396a5e7116f74c2d,
98'h35aabb2b5ff6b97fd5685d2ac,
98'h32b70ba5735781a6b983a3530,
98'h0904a8521cd4a9f9a9765492f,
98'h1fcd2e7f901d76e00bfaa957e,
98'h199d96f31a3cfd746cf6a519e,
98'h32b72aa5545043e8b1c1dba38,
98'h1eb5bafd4c514458aac1bfd58,
98'h347eec28e75d1d8e96f7026dd,
98'h024755c487f4124fe28eda052,
98'h2c79d618e361b886d3f6e3a7e,
98'h0f1b01de38aea5b171f269e3e,
98'h1d80b17b19b90ff36dce705ba,
98'h0f83b5df11ab50e3484bc1b09,
98'h09fa4f53c20bed4403018f25f,
98'h35b4912b7d8e9f3b3cd0cc19a,
98'h3612f5ac38f731b1dbc289d77,
98'h099262533b2941b6512ee9025,
98'h012a85c25d49ddfaa79d18ef4,
98'h2f52ee9e89acb2534e3fe83c7,
98'h3fb3633f414cd8c2b0400f008,
98'h222bf984523c9ee46d1a261a3,
98'h296c1b92c4767848eb78a4f6f,
98'h12c40f658a670f54e74ac7aea,
98'h010dd2421d5bc9faa79a670f3,
98'h360708ac273d500e5751162e9,
98'h3e39623c5fa198ff7776becef,
98'h127057e4cf7797dec879fbf0e,
98'h049d4bc93a1f39342faf213f5,
98'h3bcd0bb7983d6f7055029ec9f,
98'h3ffe59bfc2550cc4b094d9a12,
98'h0be79cd7e7dcdc0facf11e39e,
98'h1ffd097fffc8ccbf97f1758fd,
98'h3d7f70bae7ea450ff95a6d72b,
98'h1421b36847c9914fa6fad12e0,
98'h3a5e2434a8f31d91f8d45071a,
98'h1ce97379f48d99a9345dc348c,
98'h294c9392891d4b520c9a77b92,
98'h353dd02a558bd36b12b268e55,
98'h3119a22200bd4dc16c75bbf8e,
98'h0cf12359fe63243cd2d511e5a,
98'h36d4c22db81d29301bbc7ad76,
98'h3489c0a911916fe33186cc231,
98'h32ce3ca5a45e0c8895cb124b8,
98'h00d5e141a8ac61914a6090b4b,
98'h0ddf395baa8eb9150e1b7c9c2,
98'h3d72473ac8bdf3d1518c0ec30,
98'h2aeb8795dbc0abf7b1ab0ce36,
98'h0c9da7d902d6b745a3dd17c7b,
98'h0b7f25d6cf16045e06a54a8d3,
98'h3c62d338f2d7dba5bbceabb7a,
98'h3dd988bb9b722c76f652ed4ca,
98'h31539e229ce6f979f38ea5e72,
98'h32a8a4a545a7424b6e13f9bc3,
98'h39be873370ed95a1faab07355,
98'h1525b4ea4daa3edb68b3fcf17,
98'h35791eaad6f66dedd31be3262,
98'h0535c34a6987dd132baf68176,
98'h2a093294132a7de66f4cec1ea,
98'h3c9ff0b91b8444f716090d6c0,
98'h2526b20a689fc89113719ea6d,
98'h325b7da4b5ff6e2bda16baf41,
98'h24405788a31be10611d70e23a,
98'h156791eaf7684eaef333f8267,
98'h22dd1085b55c302a960e502c0,
98'h378ec22f3eb8bdbd7d91dffb2,
98'h1f6426fedf65fd7ecfb2891f6,
98'h13e85c67d9a41df36b631e96d,
98'h2206248432d038259535972a6,
98'h00d96cc1a4d2c489896b0c52c,
98'h0830815045e8fecbc38660070,
98'h2dc7861b903423606f7eea5f0,
98'h142605e85608e66c0a8bbb151,
98'h059f4acb21a1ac8349d03dd39,
98'h3005f7a0395602b2ba56fe94b,
98'h0cc0b3d9b2bc7fa54fdf4cdfb,
98'h01bbfdc36ca8af196b992b373,
98'h0ed3195db01fce200fbcb9df6,
98'h0602cb4c3f34163e514db8629,
98'h0b72fa56fbb2043771c93fa39,
98'h37d3852fb704782e1bb5ff576,
98'h039b85470e0eb25c046a8de8c,
98'h3b4bed36835535c6afa848bf5,
98'h311ddea237b3322f5a3444345,
98'h23454586883096504add76f5b,
98'h09682bd2fdc8123b91cc0f839,
98'h2385fe073dbb4f3b78505350a,
98'h114e5662ac113a182f57e41eb,
98'h22a8178560fdcd81d0e97941c,
98'h347699a8e1bed683758d5c0b1,
98'h127e4f64c7ed3ecfc69ae38d2,
98'h247bc588c588fdcb0a8130d4f,
98'h07f2044feae65495ccb616396,
98'h35c74babbab019355c1dd9383,
98'h2803e1901ebbd1fd51afece35,
98'h1e95027d102c0d604bb043f75,
98'h32c944a5a7eacf0fd6ad04ed5,
98'h2382af07018421c32941b4329,
98'h2af06615fd76c53ada19cad42,
98'h387d50b0e979a992f87dbe90f,
98'h1c8541f91c5f52f8ae39253c7,
98'h28ce219185df6acb8bab63174,
98'h04613e48ef91c61f2cfcc11a0,
98'h117965e2cda7c4db47c84aaf8,
98'h1edf94fda7a8640f51a1fe433,
98'h1a10ef742a639b94d11d22c23,
98'h1c207a7865b9718b50767b00e,
98'h3d8c66bb111bfee213aa19674,
98'h2e55061cb0e7f8a1d7cf3faf9,
98'h1aa9557547a08ecf689279113,
98'h073ddb4e4b585456a4a58be94,
98'h05c4e94b8714a8ce033664866,
98'h31368f227c9a75393b744116e,
98'h311180a22eb54c9d77f1b34fe,
98'h29d7d293898bebd32cd8ef99b,
98'h0f79f15ec681c44d257eed6b0,
98'h0c6a58d8f023aea04f2381de4,
98'h16748eecf4a10da952c567258,
98'h1d14817a1489a4692c678978d,
98'h0f77f45eee0e019c0f617d7eb,
98'h2edcbc1db84be9b0b9ca29739,
98'h3eb38bbd5f443c7eb77df20f0,
98'h1a4ab7f49073dbe0eaafa4f56,
98'h1e1dd77c3857c2b0b59d668b3,
98'h14a142e977acdc2f531387c62,
98'h05da75cbbd116fba30baf9617,
98'h1c5af7f88a9ede5509be75936,
98'h3169eea2e15a178294b101895,
98'h2ac3a495920eaa640f3493be6,
98'h20053880206e7200f01ceaa04,
98'h183871f07445e928b31f96c64,
98'h31f700a3ce05c1dc0fff309ff,
98'h2cc8cb1999b4e9f3719f6d434,
98'h18b4b2f167c53c0f901e7bc03,
98'h1da2077b7bb029b756548c4ca,
98'h0fe9415fd70a326e29bcdcf38,
98'h04dfcf49939b9ee7261edb8c3,
98'h1e93affd2b44f716b27629c4f,
98'h210b488210c5bce1ac744158f,
98'h2ccb561987ce89cfad2677fa5,
98'h27c2fa0fb7a43eaf77d9ce2fc,
98'h08abed515952fbf2a87fba510,
98'h1fb5777f5214aee40c728998d,
98'h1f5b53fe929a99e50c7d7b78e,
98'h1548c4ea81b2ae4365bedccb8,
98'h320b18243aabd2b57b2dbab66,
98'h3ef8843dcf45fdde938fa0871,
98'h0647bf4caaefe215ec4de858a,
98'h16a4d86d58ba43716bd7c6f7b,
98'h38d7cd31873435ce500300bff,
98'h37bc102f7e0295bc3d6fa97ae,
98'h0edc8ddda712958e2d7bc8daf,
98'h03590d4680bac2414104f3e1f,
98'h1dd69a7ba47a0d08f09429e12,
98'h0f206c5e6e48541caf5a301ec,
98'h04a0244979c293b38f98adff3,
98'h05d66ccbbcad5fb950a0f3213,
98'h315efba296e572edd2111ba41,
98'h0d5799dabb2f06b65221a8243,
98'h2ee0579dc5246e4a4d01317a0,
98'h08ce3051b561c1aaef8bfc7f2,
98'h2ac05e159e99aefd32568344b,
98'h13ae4967651d690a2e32ec9c6,
98'h312f6ca277da65afba4274948,
98'h2632c00c6a4afc14941f6f083,
98'h37171f2e29063a12180756500,
98'h22c4dc05b26e2924d54cc14a9,
98'h13d11967954d6beaaa47a1549,
98'h20e8b601e13c9482508952a10,
98'h3c918c393027be207b2e52966,
98'h11f86363e384e3070d5f519ab,
98'h091781523a2620b470cf6881a,
98'h2227da847a178034170fd6ae1,
98'h3f24e13e50791460f3e77d67d,
98'h28fb9f11f753252eb813b1102,
98'h34b03a295df5d67bf4a984295,
98'h238c26873b6723b6d7bcd28f7,
98'h03b24b474e94455d0491a4291,
98'h3ca001b96d4d6b9aba7b5b550,
98'h29e14913c30f8c462b3c35568,
98'h1ed6c3fd9cee5479cef1461dd,
98'h3e9be83d358389ab1d07dc7a0,
98'h1fceab7fa1d02303b067b3a0d,
98'h05b6234b7590f52b0ed1c61d9,
98'h0c5f0a588524564a4460d828b,
98'h0ac9c4d5a6c24a8dac6303d8d,
98'h29b16c9351f4a963cee9857dc,
98'h3a1cad342a9b7095192e07724,
98'h293383125ea1dffd51f558c3e,
98'h161edd6c24ee2109eec33f9d8,
98'h020bc7c403d64ac7817884a2e,
98'h0ef23c5dc0bd10c143ebd347c,
98'h2deae81bda7e14f4f21a3f443,
98'h205e1f809227d6e44ca17d993,
98'h14c3ece9804744c08542cc6a8,
98'h0e00955c128995e528228ad05,
98'h0f2521de649b8a892cf02b19e,
98'h197f6872cb2463d64928f3124,
98'h3d9bbd3b3af5c435fe24605c4,
98'h3eeaecbdfc637138fed3977db,
98'h10bc48e17ee546bdd3e863e7c,
98'h1c748478f7edf1afd5189d8a2,
98'h2d19c99a3600e62c38c6abf19,
98'h080ae8502674c38ccb9feaf73,
98'h24a5a689687bbd90d34859068,
98'h335e30a69b54d976b3acc2875,
98'h37a2532f5dfdb7fbf56802cad,
98'h393d9d3253d85ee793457f067,
98'h3e82b4bd25d1d48b991522522,
98'h02311ac45a10a37407106f8e1,
98'h2fc04b1f8b6c3556cecb201d9,
98'h35a08fab67f2c20ff764d46ed,
98'h34e21aa9eeb9e09d78e6fed1d,
98'h24cadf09a291090531d6fa03b,
98'h1c9e5279069c4ccd28cea7d19,
98'h213eb50242fb20c5c90e75720,
98'h3930b2b27762a62efc24d6385,
98'h3d770b3ace7ef3dcf2fd7fc5f,
98'h0dafb95b5b02da760a2ca4f45,
98'h27ad728f46b459cd4b9873172,
98'h1f5a85feb9445b329627b84c4,
98'h20e41b01c6ed7c4dc9f465d3e,
98'h3c8981b936feab2dfce20b39c,
98'h20999c810455ff48a93be6f27,
98'h1e1bcbfc10fda3e1cbc65bf77,
98'h3c887d39243aeb087830da106,
98'h1deb5c7bc50d7cca28be36518,
98'h0744794e84a551c942fa72c5f,
98'h2101ee823620952c75c8a0eba,
98'h04778d48f2a1b9a54dc651bb8,
98'h32f8aa25db70fbf6d39a69872,
98'h29f0bc13cb3e42d64d4bbfba8,
98'h351c87aa01efb543edc30f3b8,
98'h25a6988b74799128f6880a6d1,
98'h1ba17c774f43c55eaab950758,
98'h263f8b8c660c728c3312ff862,
98'h095e5f52aa0af7940cda55b9a,
98'h29a1dc936b284a16553289aa6,
98'h1b3b937667fe660ff0ce7e619,
98'h377d7baec9f43353f05c6bc0b,
98'h2bae6e17440cc1c82beecbf7e,
98'h28b186115fc2edff921d1d043,
98'h304b60a0a06c5b00f42deee86,
98'h0bdf91d7adab849b4e62c59cb,
98'h1ba8de775716e96e2caff1f96,
98'h176eb26ed45eb5688af359f5d,
98'h107d0560d211126408a385f13,
98'h05b042cb43c31847825cd6c4b,
98'h3c1007b8304fb2a0bb17ee963,
98'h2cc86d99b712092e18f69db1e,
98'h09cd51d397fce76fe8728e50e,
98'h3d6c73bae4df4e89b892f0912,
98'h1bed73f7df4ed2feaecf11bda,
98'h0d78b55adfa582ff4b478e168,
98'h39e2c7b3e612278c17fd3bcff,
98'h09d079d3ab2139966d3c6cda8,
98'h0062dbc0ef7a6f1eebf752b7f,
98'h19e976f3d0f4eb61eab798957,
98'h3c9697b901ba10c34f942a1f1,
98'h02d51945afbf9a1f6ca52cd94,
98'h082b285063541c06aadfd115c,
98'h2b898e1727003b0e34a272495,
98'h22ada3057909cf3216eddc8dd,
98'h249c88090bcfe057ac1b1a183,
98'h31cb72a3a6b5df0d7620546c4,
98'h3e91c93d0aac9c55724f9964a,
98'h31c17aa3a557800ab5c63eab9,
98'h274f6a8ead3f2d9a5523a60a3,
98'h3d74033adcff2d79d69ccc2d2,
98'h3539e4aa743566a85a5bd2d4a,
98'h1e595f7cb63f302c552623ea3,
98'h10e9d661c0fb53c1c4794a88e,
98'h139154672031eb004cf0cfd9d,
98'h115d8de2b54d23aa91aaac634,
98'h213342027217dd2414d2c7c99,
98'h35f84fabe34bd286b651088ca,
98'h090d0d5235ff6dabcfc31ebf7,
98'h3191612333ee8ca7d95ffb72b,
98'h38bcc43148d8735190654de0b,
98'h0e44cc5cb75adbae9167ea02c,
98'h0a3f08546fc57a9fae8120bd0,
98'h0ea7ebdd6edd8a1d8f615d7eb,
98'h17bc366f466cd04cc78a41af0,
98'h3273b0a4f6ee4fadda588014a,
98'h258e4e0b1a7b46f4d002653ff,
98'h26a6ab0d54d835e98edfb83db,
98'h322999a4617ac002f4e91669d,
98'h0790d24f3b50c03690b864a16,
98'h1ec2177d938e76670c9423792,
98'h322b0ba46777d78ed668b8ccc,
98'h09379f52539700e70733a80e5,
98'h0d8c755b306a6e20cf7db8def,
98'h2402cd8807b01ecf6aecbb15e,
98'h313f6b2252c1e96591005521f,
98'h078ca84f17ea3eefe7ddb9cfc,
98'h35a84fab530a49e6122ca6645,
98'h2d8b091b1091c5610f87339f0,
98'h0ca015d9526913e4e7c24a6f9,
98'h2eabc51d5d46177a92fc7725f,
98'h15d485eb8b5ef4d6a84cdeb09,
98'h010893c216925eed05e6bcabc,
98'h387048b0edbe2f9b598b9e130,
98'h068db74d28aa16916bcdf377a,
98'h3dfcad3be49fc00918a71b513,
98'h01ad65c34b5b5056a3422d868,
98'h355f312a83514646ae2c1ddc5,
98'h3069efa0d538bb6a5168aac2c,
98'h2444ca0892e5ace5edca9dbba,
98'h25f0a88bc26d6ec4ca1785d42,
98'h3d3cec3a4d4290da929fdf453,
98'h2daf8f1b4e9c70dd0f12fffe1,
98'h0d36525a68346b104d5aaf5aa,
98'h1bffb577dc9dfef92e276d1c4,
98'h17ff866ff74377ae93d0bf879,
98'h1c2e677852dc9565abc2bf378,
98'h04dd29c989b35cd343a421a73,
98'h15df146bab83b6171058b2a0a,
98'h0637fd4c4f47945e855fe46ab,
98'h186ff7f0f8a274b154449b288,
98'h2dd4a69ba616928c34face49f,
98'h263b7f0c61d3b9039203ce03f,
98'h1df73d7bc9e5afd3c9f73b53e,
98'h2740730ea6ee4c8dd38bafe71,
98'h1b448df69e37ce7c6e5f171cc,
98'h06eadecdd5ae9d6b47265f0e4,
98'h2723238e4368c346caa2f9b54,
98'h3767b92edb3c4a7654a900e94,
98'h1ace137580df7f4186eb64adc,
98'h121d4c6409dd67d386fead0de,
98'h343b7e285690f6ed32b31d456,
98'h3c925bb90b1989d631eaf963d,
98'h0368dd46eabdc7954b89a9370,
98'h273e100e62fe8c85f28f27251,
98'h248f08891204a4642da4eb3b5,
98'h146a9b68de29197c6ca4ed395,
98'h0e2fffdc4b9378d72670de2ce,
98'h2484a3891da2f17b7089e5412,
98'h2ce07099c57154cacc9471592,
98'h16e1696ded98f51b311e97a24,
98'h2e1f001c018b12c32bea84b7d,
98'h0e35afdc4a5aeb54862426cc3,
98'h337b52a6cf5cc05eb0b604c16,
98'h22a7660566070a0c322b9c046,
98'h0bbed3d76bc1c697ade0269bc,
98'h2c940d9904b33f494c51d3389,
98'h3cb93cb944a5d1495057c380a,
98'h26d5e38d98d635f1afeb065fd,
98'h39c2df33850075ca0fb0d53f6,
98'h1981c6f30a2221d448e8fa31d,
98'h14f6ab69fab59f3553eb12a7c,
98'h1ac7e1f5b9f344b3d52ec9aa5,
98'h2795f78f07a4b14f4bceaa379,
98'h26d1130d85e438cbcb2d52f65,
98'h14f80ae9ed60741ad0961fc12,
98'h052312ca7709f4ae0f0b41de1,
98'h06d761cd8bb9ba5744a447093,
98'h36455c2c96c9986d9343bd268,
98'h0dbeb8db6976c892cdcd605b8,
98'h2310d6060529f14a4a0eb1d41,
98'h08c7d351804180c0a24255049,
98'h0c443ad883f2c5c7c40dc0281,
98'h18ce02719506466a2b751236f,
98'h30a73e2171dbd8a3b8a0c5b14,
98'h08a6705150ada6e1465505cca,
98'h1636786c457db64ac6ed0badc,
98'h39e02433de4ac57c960aba6c1,
98'h03820b4734a637a94e0a10bc1,
98'h27fdce0ff7887d2f17e192cfb,
98'h0d990d5b3622ceac70eef701e,
98'h2f0b4b9e0a4f4ed48e56a69ca,
98'h188baef12e028a9c11a38e634,
98'h11e0f263ef4e049e904bbdc09,
98'h10be236172c1e3a590e001c1b,
98'h3c5695b88c3f1c5872256c844,
98'h25f6490bf0c23fa1b5ae222b6,
98'h0a1851542274ee04eb234fd64,
98'h3a3e12b45cdf3b79b5c7538b8,
98'h2fbf0f1f7e66963cdb8969570,
98'h3264ac24e2e3b285f55217aab,
98'h1d3ed07a6ba79b1752399ae46,
98'h301864a02510890a354a3b6a9,
98'h0aacb4d545e4564be42442c85,
98'h22435784b2d73125b546a22a9,
98'h36cec42da72d1b8e577ef7eef,
98'h1384d2e73259f3a49177b1a2e,
98'h2dd7741b9a0a247431f86623f,
98'h1c517e788e33f85c4aa15db53,
98'h121ef1e40682324d2628490c5,
98'h2a744514eb7b0e96d57bd4eae,
98'h149c29e9186dfaf0eb4289368,
98'h1659ff6cb6dd34adb34dcd069,
98'h2b4f8e9687224e4e6c9c77394,
98'h0bc1d5d7972bdfee48bb6d717,
98'h1cc1a2f9beab013d76db290dc,
98'h0b1c6cd6039703c703acdc274,
98'h05273f4a5d80927b08a9f4715,
98'h0713ccce3849dbb08fd76a1fa,
98'h07ad9c4f52d291e5a6a00b8d4,
98'h0a660754c90b725204dc5e69b,
98'h08e018d1d530cdea478439af0,
98'h316ca322faf4e7b5db1862b62,
98'h1209c364338d35271165be22c,
98'h045ac048983f7cf047268f4e3,
98'h34e4a0a9d74082eeb30948e62,
98'h2f6c029ef79c58af19c216d37,
98'h2ed8b49db8eba3b1f9f11613e,
98'h20ee3801ef78111ed41992482,
98'h3f7ccb3ef7bfe1af5dcf2b3b8,
98'h063fc3cc40fbf341e1ceedc39,
98'h22fafd85fee7c7bdd878b150e,
98'h248cc0892a8f0b9513c6f3078,
98'h026afd44db7acc76e779726ef,
98'h2c44ef18a208ed04139377072,
98'h2e241a9c6295b885142e74c85,
98'h12f45a65efb8399f70ab25015,
98'h34790ca8f6e1d2addad6b7d5a,
98'h0258bec4a0ceea81a8c9ea519,
98'h1e3f79fc6b04c09612510ea49,
98'h313db5a245b6584b4dbd037b6,
98'h25f53e0bd723366e4f461d1e8,
98'h0ed99add8b3d01564685a70cf,
98'h1a4576f486d0584da84573d09,
98'h38153430308014211a2552144,
98'h251f460a1673e86ccee4cb9db,
98'h03581c4682e2b5c5e18eb4832,
98'h21805f03376128aed63861ec7,
98'h3723e72e61550a82961e3c6c3,
98'h1f854aff0c8889590b0375160,
98'h05f80ccbec9cfd190ca542793,
98'h2c417018b2de0aa597c7deaf8,
98'h1aa88ff57742c8aeb47ad6290,
98'h0550dfcabc3e6a387063d280c,
98'h2781648f19333cf2702d28606,
98'h0b05d6d635cd072bb034b7807,
98'h34409da8bd19caba3c569a18b,
98'h23840a872f748c9ef4be25c98,
98'h1f214dfe6be44917d2c165c58,
98'h110bafe22d64579acf9c01df3,
98'h17e1336fc1d27e43a66cec6ce,
98'h1a2640f46214a1042f0eb87e2,
98'h14db2069b3e367a7f22fa2046,
98'h075707ce938b64e706b89b2d6,
98'h0e00215c186240f0c99898933,
98'h036166c6cd4c095aa42b5c086,
98'h33a965275dc54cfbb45bac88c,
98'h1526dcea458bc7cb26aca92d6,
98'h0bece857fc005e3811fb51a3f,
98'h108ed16113f4d567e920e9b24,
98'h2c4ed61891dd1de38f8afcff0,
98'h3ada1ab58e72495cf2531904a,
98'h1359b96685db144ba64d336c9,
98'h12344664412ec64264d8c329b,
98'h01d75bc384897049019833032,
98'h2c449f988e1fe25c2e99207d3,
98'h0a147554113c8fe266d4414da,
98'h0ff0fa5ffa284db4728652051,
98'h28c90f11ad71481af58e95cb2,
98'h077437ced60abbec075fbceeb,
98'h0aefadd5db1fedf62983e6f30,
98'h055a91cab4178c280e5c877ca,
98'h320539240ab11b554f2d951e5,
98'h14e5a069c4af2f49666533ecd,
98'h20dba3819a363af44ec4779d7,
98'h08ca2251af63529ece0b5d3c1,
98'h2a59529484f7ce49ebd44837a,
98'h2e29861c58b0c5f171b693037,
98'h0d2f475a7c5b74b89262af04b,
98'h111930e228fc2291ce8554dcf,
98'h07c0054fb993b5b33054eec0b,
98'h17f986efe4ab37896f292f9e5,
98'h2a213a14667b878cf42730685,
98'h3f4eb23ea2e52c85d88cf7b11,
98'h2d52291a9f6f97fed33070465,
98'h0cbd2e597cb36e39725c2724b,
98'h2a70cd94c3e751c7eb9607d73,
98'h013c0bc254ed5269c58a578b0,
98'h3ee7c7bdebffa817fab9dbf57,
98'h247efa88e688820d12c1df257,
98'h273f020e62199e8432562824a,
98'h120a1264069823cd26288d8c5,
98'h2d691a1acd1e8d5a2ea1e9dd4,
98'h3751582e8574bd4aef31855e6,
98'h1d1788fa05ec2c4be8c0ed518,
98'h0db60a5b4336e246643b3b287,
98'h14cf8969bcda5ab9b46a7908d,
98'h0723a4ce6ade9795ac808f190,
98'h2929c212573ca76e50199a602,
98'h3c7ea9b8c9317f52716c0a42d,
98'h34d6ada9a4319608564210ec7,
98'h2e072c1c2489bb0914a439c94,
98'h07b1c04f7001ac200decdb1bd,
98'h2b411496857f9b4aec302bf86,
98'h3d5d513ab1c034a39bc761778,
98'h3de42c3bd188006333db0b27c,
98'h049143c90bcfc957a41843483,
98'h15c5e0eb9c518778ac85da191,
98'h17766ceef95c9b32b434c2086,
98'h2e9ed19d36da6fad995e5052a,
98'h3f18bcbe04ce7ac9b0f9cde1f,
98'h17fe136fefe9449fd1f9d603e,
98'h042a284861a49e836973b1b2f,
98'h27ac390f7cc24339991b9f123,
98'h12004d643b1d2d3633475ea69,
98'h0b30205646a3844d6474e928f,
98'h19e6ddf3d47a83e8eb9858773,
98'h221770842dc1e31bb3f654e7f,
98'h2090c60133a83e27550e410a1,
98'h2414ec882130a702515164e29,
98'h19a216735772006eec4505b89,
98'h0ff674dfc04de940841117881,
98'h39fca833eb6dfb16d95aa8d2a,
98'h16e4ceedc1fdbe43e638a34c7,
98'h04a989c9612d38024975b072e,
98'h264f318ca42e1d88529f53c53,
98'h33e92427cc33a058700731201,
98'h36548aac96cd8a6d934885468,
98'h0c2422d870a9c1216f3378fe7,
98'h166c856cfc8e79b934bebfc98,
98'h0d271b5a5faa5a7f6b345d767,
98'h3282552525817c8b1600f46c0,
98'h2342f8869b7da076efb0263f6,
98'h33a33c275fc026ff94d8d8c9b,
98'h199c1ef30e04475c29e81993d,
98'h0cd2d4598d12b65a067962ace,
98'h2d22559a78044a303949a7f2a,
98'h3287142525aa7d0b760c644c2,
98'h285b6f90a4f97389d35538c69,
98'h05be1bcb5bbb07f7485e48f0a,
98'h2f5ab21eb87ba430f9f59593e,
98'h1e8fb8fd3dec063bd71eefce3,
98'h04eefe49d43cdc68664af6ac9,
98'h398cb1332b4df2969936a8f26,
98'h2241b784bc1103383794aeaf3,
98'h132dc86676ab7b2d727650e4f,
98'h24d06c09bc616eb8d84c76b09,
98'h110489e224c1a789ad718c5af,
98'h27db3e8f8ade2c55acae5ab95,
98'h354fcf2a8d18c4da309a25013,
98'h02120ac41d2f077a47d0448f9,
98'h1b060a763be80837d5bb84ab7,
98'h227a5004e1d65383911428e21,
98'h1a574a74909dfbe12abd51957,
98'h1437da6860677300cd27d35a4,
98'h141907682457a488ae1c2afc3,
98'h141225e823a31f076ded513be,
98'h397da732d1c069e392cf84459,
98'h08408bd0adfb6f9bed8efedb2,
98'h10e9c6e1f084be21305ba140c,
98'h1f3727fe7371a426d4aa33094,
98'h34a9422945b187cb4e96b27d2,
98'h08de80d1a6afa98d6be38a97c,
98'h30b5fca17c0a46383b3010b66,
98'h32cfefa5aeaf669d785fd590c,
98'h35b268ab778ffdaf3b509996a,
98'h17e0c96fd231be644a84a1f50,
98'h2ca9cf197222dd2457b32b0f6,
98'h197645f2eab75c15510b68820,
98'h0d1857da1058a5e0a75c3f6eb,
98'h29cc2793bd9d3a3b39da5873b,
98'h092cd2527151d422ae9fa99d4,
98'h1588246b0b6ee9d6e83dc3908,
98'h2f263c1e6e87889d376b712ee,
98'h24a40b8977709a2ef705296e1,
98'h1e1f0b7c3d3c2cba56d6ce0d9,
98'h22e8b285f7d2e3af96aee58d5,
98'h1c8833793668deacf4bc44898,
98'h12e397e5c5f24c4be635790c7,
98'h1b05ef761fb1977f4eade1bd5,
98'h27714b0ee1749002d23976c46,
98'h335049a6b41a11a839da96d3b,
98'h0ba69b576505ac0a0c2b11d85,
98'h1c29637849e57553c983b6330,
98'h0b1276d603e6a347e3be46878,
98'h156b7c6ad83abaf06b698dd6d,
98'h01029842087007d0e25ca804c,
98'h15a0bc6b76d7d72db31e24e64,
98'h20a4ed01711a42a2346fcbe8e,
98'h0186b8c3084da250827516c4e,
98'h158fbf6b0f8d9bdf294756d29,
98'h094fbed2bfee7e3ff24f8f44a,
98'h386a9930efac029f5a05a6f40,
98'h2b63db16ebc9c117b5cb670ba,
98'h0a21f1d44776954ec46621c8c,
98'h2cd3a09984bddbc94c645f18b,
98'h253f920a6020e88071581ea2b,
98'h109eb1610edb415da7de7cafb,
98'h04b1c04948941151035174669,
98'h14600668f702102e32d885a5c,
98'h2d7b221ace1369dc2ee3a2fdc,
98'h36e1f7ade3d47a87b6ad9c8d6,
98'h21756b82eca51c997386a2071,
98'h278c048f0bc7ecd78cd4fc59a,
98'h1080c1e102506ac4a4b44b297,
98'h308c5ba11c4ef6f89336d4a66,
98'h2f29e59e4a33b4544e57667ca,
98'h150f216a02c5f2c5a5f5450bf,
98'h3a011a341ae440f5d53956ca7,
98'h34c57a2982fc6ec5edf07a3be,
98'h278bce8f1279c5e4ce81651cf,
98'h2a6e5094e4e55289d3d4e8c7a,
98'h2beb0417de17b07c3280ad250,
98'h0802e0502f27cb1e6dcaaadba,
98'h2500778a1eb62d7d50eda941d,
98'h2498f8090afaee55ebe4f997c,
98'h180c88f02d5cef1a915a5e02a,
98'h21fd0a03dae625f5ef38cbfe7,
98'h066ee24ce9f1b813ec1826983,
98'h3e75ecbcedb0559b7b0990961,
98'h1263e164ed2ca19a6fe420bfd,
98'h2e14659c14f7c669f0c30b018,
98'h2248be84a4342388519f38833,
98'h32607324ef9cca1f387f4f510,
98'h3520762a66d2dd0db6fcd4ce0,
98'h332650267759272eba9fddd54,
98'h19c36ef3bc291cb8557b22eaf,
98'h13954067028e3d452588df6b1,
98'h3f53e13e992c26f27620020c4,
98'h1fd215ffbb83f03736d5818db,
98'h0d4102daac3540186e5d90bcc,
98'h148f796939024f3213647226c,
98'h2752ea8e9d52737a912957824,
98'h282df390755ffb2ab7637baec,
98'h22e93b85c7fb1acfcab915956,
98'h3f55b3be84cf5149910941420,
98'h09c68bd3b43a27a86f802cdf0,
98'h11ec1763ede4511bcff41a1fe,
98'h00728b40f7502a2e8df0ad5bd,
98'h14b6f3e953fd44e7ea2d0e345,
98'h0e6ced5cc23f1944642b01a85,
98'h3bef9d37c6682a4cd095f1e12,
98'h091b11d23ba1dab7512f3b225,
98'h3777aeaeecceda19b911a2322,
98'h0b8a68d72da18c1b6e4afd3ca,
98'h1e51927cbda3f0bb56fd60cdf,
98'h20d1a0018cca8a59ab670a96d,
98'h386ec9b0d9fa7373f49a4f493,
98'h210a870204f336c9c97f6f72f,
98'h2fd5f41f9f623c7ef3ce0c27a,
98'h258eb80b0a5684d4abf94f37f,
98'h08929951281320102c296e585,
98'h3451012882743cc4cdb14f7b5,
98'h0dd0af5b97e0d6efe96c6192e,
98'h3fdd8a3fae39079c7b85a4770,
98'h05f5e34be521a20a4ac5e1558,
98'h25babf8b71603422f5c6bceb9,
98'h337aa126d3e1b8e7f1d71683b,
98'h1b94f7f71df1407bce618e1cb,
98'h08b4dbd1436d6ac6c30891a60,
98'h08cedbd1aa2b21144cbe7f397,
98'h3db6963b466c0bccd108a8820,
98'h09c09153a71f4b0e0c37f7186,
98'h04d228c9b0759a20cd51f0ba9,
98'h181f9ef00aae795568b386116,
98'h28464b909d3d287a7160dd02c,
98'h3cb997b9648935093850b330a,
98'h0603de4c211a020229c778139,
98'h0ddb815bbf4620be934868868,
98'h216f6e82dce99779cf96417f2,
98'h3f6ffcbef88ffc313dfffe3c0,
98'h3a7081b4c3f422c7ef99291f3,
98'h3a0e2cb421dd6d83b6fae68df,
98'h01109bc20dae125b43afab875,
98'h38e360b1fa148c343cbdfb398,
98'h315c0822bae02e35db0f0d961,
98'h1f9179ff23ec2487d0df67a1b,
98'h2026608051f081e3ec85b8991,
98'h3ccc14b9a0ccc281976635cec,
98'h22c4d685acb6041973deb6a7c,
98'h10ae716168637a10ee447adc9,
98'h3dc03a3baf70ff1efb4c4e56a,
98'h1a741a74ee086d1c121f21e43,
98'h04f0c249f03236a06d48be3a9,
98'h346e4ca8e28b140535be582b8,
98'h0e6594dcc42ad34864a41a095,
98'h0ac021d5bee647bdd2699a64d,
98'h24ea0f09c10f0642097e4552f,
98'h0d9b74db3ece06bdb31a5ee63,
98'h02eacdc5cfe576dfe4b411297,
98'h0e688cdce4f8ff89ccd86319a,
98'h26ec738de04d640091ce75e39,
98'h0c7282d8ca77d754c5ba968b6,
98'h03b632c76b759296cbcaf1578,
98'h3d626bbad25c31e493efa767d,
98'h03c213c7b0adf1214d1c013a3,
98'h24033f083f617abef8d92e71c,
98'h0d74ffdaf6ae00ad5108c0220,
98'h38787fb0d6396bec73ac7ae75,
98'h081084d01059fee0a61aa0ec3,
98'h0c41a358888e56512533fe6a7,
98'h0c4061d8b600c9ac30904ae13,
98'h1e143a7c16bd2a6d4d34593a5,
98'h0a95cbd520bc8c814ad496159,
98'h09c6d85384b93ec963a005c74,
98'h023276c448d0265182c0a7457,
98'h1336bbe6657bd98aee2ca55c5,
98'h3e555dbc9d8b4dfb16f82aede,
98'h044236c8bbd178b7b004ebe01,
98'h366b4b2cd16f7f62d1f6b2a3e,
98'h21a1d5037b46d7b6973a2b2e7,
98'h35b51fab53ffa167f26d3044d,
98'h249a47892c67ba18d44080687,
98'h1985dbf317d46def8c569278a,
98'h1c31087858717170cd289e7a4,
98'h1b8a66f73b3f993675b2800b6,
98'h23bdc487460b274c0a723af4d,
98'h3c7d1638dff7bb7ff71d346e3,
98'h2a628514f685e32d383a1a108,
98'h1716f7ee1ef6f67ded837b9b0,
98'h232496065596556b0e2ebadc5,
98'h2700d68e1ce66079d0f9cdc1f,
98'h0c102dd8286a5a90ed1ea21a4,
98'h3ff6073ffd2029ba7f458c3e9,
98'h1800d570186c4970cc1b47b83,
98'h0a3aead45982867308ef5c51d,
98'h1658926cb5f5f4abf313a1c62,
98'h36f93aade7fd540ff7bda3af7,
98'h021fcb441ba57877677150eee,
98'h3d040f3a1ff485ffd73e254e7,
98'h1ab7f3f56ff5be1fd2ab6c854,
98'h28f5a791ed41471ab58dbbab2,
98'h177af16efc2cc73854e9ee29c,
98'h1e88f17d18cbe7f1add5365bb,
98'h195143f2a9a1b39350bcbde17,
98'h3080d221336882a6d8fa5531f,
98'h3d78ef3acccc8b5992915ea51,
98'h2c5f2d988ad065d58dcbe4db8,
98'h0f6722def481c32930fa39820,
98'h3b9dafb72e42391cba77fa34f,
98'h18de9f71972b88ee4c028a17f,
98'h090a51d21482e86927634e8ed,
98'h2304e1862bc2c897b3b1ea877,
98'h0a59a554bba94a377180bbe30,
98'h2d700a1adcb9f5f9528a80050,
98'h1ff0d9ffe84e8890b20fd8a42,
98'h1cd782798bfb91d7ea34c5146,
98'h0b598756a96d4792ed31b3ba6,
98'h3641682cac8e761938b3f7917,
98'h03c133c784698fc8c20ab0e41,
98'h1136b4e24461db48c566240ac,
98'h0b569bd6956b726ac83083905,
98'h0fb8235f53331fe648bad0d16,
98'h1446bbe88f66765ee8eb4c91e,
98'h095ddad29e6f527ce9f34b53e,
98'h1c8b96f908d7bb518958d492a,
98'h3c3bd438596277f2f567930ad,
98'h28aebf117274e5a4d6c8e92d8,
98'h2dd5049b88f693d1edb2e61b6,
98'h0b119e561fb5c37f4ab1d8755,
98'h3c9743b936b4722d5cd2ed799,
98'h2b3d7b167a52b6b4b9640c72c,
98'h2309f38603a82cc769ac88136,
98'h232d46067d81dbbb382bc8706,
98'h25096a8a0d3b745a6c9137b92,
98'h03731cc6f7ecf22feed803bdb,
98'h39191932180799f034482cc89,
98'h3e8b943d000a05400fa5665f4,
98'h080672d0331153a62ec5f19d9,
98'h1ba0c0f749b0d1d3495464b2a,
98'h3fc695bfbcd048b9bf25b79e5,
98'h3d6efd3ad176f0e2d3b97b876,
98'h3fa8b43f7ed4553dbf9f425f4,
98'h3eed743de68cbd8d395e8c72c,
98'h3fa73a3f70ca95a1bc1c73f84,
98'h00cc6641aa84ff150ad45955a,
98'h0ed1b85dbc142d3812b979656,
98'h3ccb33b9b3a14f275c1b20b83,
98'h09798852ca10ce5424e295a9c,
98'h2a58241485ed424bec1159982,
98'h02fb3845dcaf01f967ea8e8fd,
98'h2edbed1d9da24ffb531f8f463,
98'h3caeb03966c42f0d98dcb7d1b,
98'h1782fbef35fe7aabf3605da6c,
98'h2fb81c9f6c1e669836f5a0cde,
98'h2e467c9c9ee7b7fdd34b8d269,
98'h162393ec5c31e5f84c955e792,
98'h3c6722b8fd6618bade734edce,
98'h0ce57f59f9b461b351a678434,
98'h357bafaacb2eb0d6702a98205,
98'h0809c35031680ea2ee5c747cc,
98'h33a53d277c293e385bf39ed7e,
98'h308ba7a11ec867fdb3d503e7b,
98'h1b6b4376ea0a9314315d75a2c,
98'h0c007fd8223ab6844b8ecd971,
98'h083160d071cdbc23ae7fc73d0,
98'h0d6f10daf5d45dabb0d0dba1a,
98'h0528e44a5905e872078bb32f1,
98'h105dbae097b8dbef6a05a5b40,
98'h2e10121c05b3134b4cf0c959d,
98'h0f5161de8781984f25b4be8b7,
98'h1b012ff61e73697cce5d265cb,
98'h11a714e3731169a6312e1fa26,
98'h0f0346de369b742d3167aec2d,
98'h1de274fbe2a5dd05502214804,
98'h3dfeb23bc5eefecbf0fb6c41f,
98'h213ade8277e83eaff648c74c9,
98'h002763404264c044c0a308e14,
98'h3f6152bec430614870e46d01d,
98'h2adee9958f8ec25f0e9b6afd2,
98'h0a291a54531b26e60751104e9,
98'h25803c8b06f188cdeb1c71564,
98'h03ed33c7e406c88809fcff13f,
98'h2777420eeac3fc15948ecf891,
98'h353c77aa6af6df15f80cd5b01,
98'h387617b0cd420edab16e09a2e,
98'h128682652bd22917af962adf3,
98'h078a19cf25ec258bcb5d8fd6b,
98'h1d3358fa55dc156bacc3db998,
98'h1642aa6c9fbd427f4d7ffb3af,
98'h20bfd5814cbc07d94b5ef756a,
98'h060bbc4c2b91e8172c676918d,
98'h1428cde8445465c8861f4cec3,
98'h2b4e1816bca9c53979fdf7540,
98'h0e1ef85c191b597209ce94738,
98'h1fd7677f965e1c6c8d8d60fb0,
98'h0b2d97d65b975d7709b13d535,
98'h007bf7c0e5d6e88b8994b8131,
98'h0c2de258771182ae30cfd941a,
98'h0cd447d994b8cae9486344b0b,
98'h3d11283a2d7f799afaa428754,
98'h1f684cfefe75ad3cd7777e8ee,
98'h2c3bbd18711759221754c58e9,
98'h248a7a89051a2d4a2a6929f4d,
98'h0d5a9fdaaaef2715ce1271bc1,
98'h32948ca51821c3f052ad94255,
98'h1bcde1f7997a2172ed5200daa,
98'h2b280c96640bac0813ccee279,
98'h1c71cff8dda5c3fb6e85e4fd1,
98'h36849c2d001a8d400da7ca5b4,
98'h08c0d8d1a5c8908b8ba25a574,
98'h33f5fba7d4d8e0e99233b7245,
98'h01f83843e6849b0d0a1f34d43,
98'h00cbd1418dac1b5b439dfb273,
98'h16195bec172fcbee6b5249f6a,
98'h363d33ac7df0943bdd0b71fa0,
98'h0e520bdcad43eb1aaee57dbdd,
98'h1209f06422c82e85ad3487ba7,
98'h3a85533534c867a9bbd36eb7b,
98'h219b920321f5bf83d0e45461b,
98'h245f29889e97e0fd10bdc2a16,
98'h17d82defbfcf37bfb5e9d96bd,
98'h118cd8e30cd36a59a79810cf3,
98'h2ec8e49d8e808b5d0f525bfea,
98'h2c642418c5c5984bac8a6f192,
98'h33a62fa77b8958373bcbe1f7a,
98'h187334f0e1e74703ce969efd2,
98'h19cbe773a98f509330d6ce01b,
98'h11233be27ea81fbd53f2d6e7e,
98'h0b870a57204f6100aaf59ad5f,
98'h3fc7e03f990ce3f21635310c6,
98'h229f470516a7996d4e51b81c9,
98'h282561906d25739a7552b54ab,
98'h19ee42f3df63d37eee54859cb,
98'h2aa784156dcc959bb61d066c4,
98'h2146a1029ca71cf96f7b6f7f0,
98'h163336ec571380ee2b51adf6a,
98'h215cce02bb7bdf36f7362b4e6,
98'h24acfa09612b2182517606e2e,
98'h2a538314a544c58a93e61227c,
98'h30fe0c21ed8d241b17a2cc0f3,
98'h18fe11f1fb786636d51d9e0a2,
98'h07924b4f0896bc51040a41e80,
98'h30da69a19f41abfe940705680,
98'h0ef8e25dc2b72b45446c0368c,
98'h1734e26e664ef98c8f60f6feb,
98'h3981afb311c40b6392d16ec5a,
98'h02d7c145bc4a18b88fc8767f8,
98'h26616b0cd8f55371efd5af9fb,
98'h2f18841e3922dab25a0ed7b41,
98'h1d1690fa007b22c0e7646ceec,
98'h2d04e71a338685271822db104,
98'h0c7906d8e88f47910d42139a7,
98'h25e1ad8bf88df931179be9af3,
98'h3c0e87381b54887695d8c3eba,
98'h031d28c621dc9a83893e70d26,
98'h15edc6ebe8c5a7118facdb7f5,
98'h154782eaae19f71c10d85e81a,
98'h25aa5c8b6c663098f48423491,
98'h3992c2b310e031e1f29cbd254,
98'h09736bd2d956fe72a8b29a916,
98'h3fcc98bf92e925e5d4ad6fa95,
98'h29bf09936ae08115f527e2aa5,
98'h2db3e21b5d74537af2ca0d659,
98'h058c674b3974c932efc04c1f8,
98'h0bfbf4d7d88f85710922de923,
98'h0976b7d2d29b4e650704818df,
98'h293fa412671c388e3416f7282,
98'h2a82d995092876524cead3f9d,
98'h0b960bd7311bc6a20f2c749e4,
98'h26c1bf0d9e92ddfd11552742a,
98'h1e6b15fce0fc4a81cfd9d81fa,
98'h099194d3222861044aee7d75d,
98'h23adc28767504b8e92bf83857,
98'h2b77a916cb54e3d68db3233b5,
98'h095633528d8b22db25b8558b7,
98'h0a3d1854651cd78a2bd67bf7a,
98'h1ab56ef5480c245008b064d15,
98'h11282f62765d862c91e16d63b,
98'h13f0eae7ddf288fbec78dcf8f,
98'h26dc968da8551690b3cc6b479,
98'h017bd442cde412dbe3d7f9c7b,
98'h229c39851f64597ef08024c10,
98'h095018529e20777c69dc23f3c,
98'h1152efe284ec4b49e58fcecb2,
98'h1c1929782feb869ff3012c060,
98'h0006e24000996241002811204,
98'h1572896ac68815cd26fea7ce0,
98'h00f7b541cf5e925ea41591e82,
98'h1fcc11ffa4ada289511e6d223,
98'h1ee6717de2d21605b06e21e0e,
98'h3e75fabcfc92be391ec22e3d7,
98'h1ab027f5788df8b134cf8829a,
98'h0ac6a3559a563674894736728,
98'h2e955f9d02a65a454c4eee789,
98'h343c19a87ac0f9b59bbf44d77,
98'h143838e844377b48461bed0c2,
98'h0aeb6355d50ac36a27fd89b00,
98'h3a8b57350b7d8356f18236a30,
98'h037f8346c97b8052e33ec0e67,
98'h239b888731d807a3b55ce40ab,
98'h187a45f0d4737a68eb3b70167,
98'h134e30669d8b55fb0c3661986,
98'h2958c412a1943c0312bb40056,
98'h3bde6937a5017a0a1837f8d06,
98'h19adaff351743ce2eac87b359,
98'h3712f3ae03bd07c76eb3fedd6,
98'h3433592841774542cd6aa79ac,
98'h07d6dacf8a1fa054247d9ec8f,
98'h1447776895159b6a2a5744b4b,
98'h230edb062e963d1d34694608d,
98'h0f32b05e6e0be51c2f4fa55ea,
98'h04358e4864ad36894a38b1346,
98'h220de084199dd6f32eeaedddd,
98'h26784f0cf8fe0bb1f7dd96afb,
98'h0507254a084594d0a3532e86b,
98'h09bee4d363d8ea87ab65f3d6c,
98'h0d38a0da56d9e0ed8904a071f,
98'h0037e8c06bfbf817cb0cf8360,
98'h373305ae5064fd60f1e600c3d,
98'h08b3efd14a9a595504d392499,
98'h29cddd138a9659d52d190dba3,
98'h00497140a664f78ce9ab9a336,
98'h36bf8ead5fe8f77fd5aa218b4,
98'h266b700ce8370f1053a89fc74,
98'h30ef2a21fe4892bc9bcdef379,
98'h15cce16bbd786f3af4d15429a,
98'h1b61ed76d32f8be64ba45e574,
98'h1e1ad67c0e37895c6b1497f62,
98'h13168d663ae78d35d37f86a6f,
98'h22c762059b6d33f6cf8d257f1,
98'h26103e0c0bc6f457ac75cc98f,
98'h35cf43aba0cc3481b5a6de0b5,
98'h26437b0c8bf4f9d7cc8e1d391,
98'h1e944cfd10ee8a61cbe0b5d7b,
98'h2c068e18246e9908f41d49c84,
98'h089689d10ea26f5d45ce3e4b9,
98'h0517d94a22b6398569f384b3e,
98'h000629c03e89273d0fa3d43f4,
98'h373bdb2e5fc8147f95c0fbeb7,
98'h16d828edad29849a71006b620,
98'h23e4fb87da9d5df50fa0965f3,
98'h1837b2f06b08301630cff8c1a,
98'h394711328ab82dd550ffcfc1f,
98'h3dde51bba647b28cb90981121,
98'h10a8a8e14fe226dfe822b3f05,
98'h370cd02e0bc23ad790b3c2c16,
98'h1db40e7b7b77deb6f64afb4c9,
98'h278ee58f147f2668ef0382fe0,
98'h02fa14c5e94b0612ab1146b62,
98'h22639b84f3d64aa7958e798b1,
98'h38c89e318655504c8fc77b9f8,
98'h335476269a82fc753375dca6f,
98'h10e6e461e6261c8c4dc3403b8,
98'h18f55df1cf58d5de8a138cf41,
98'h3fb97ebf7124dba27c3796987,
98'h09374452733c41266f1ce15e3,
98'h0dc02cdbb1723b22cfcc99ff9,
98'h09e78f53ff70c0bed2561404a,
98'h274f5c8e9e620a7cf16c59c2e,
98'h38263fb0673ef30e77d94cafb,
98'h07d7734fab37e3166cc3d5998,
98'h1a0cd9f41c646078ed9c4e9b4,
98'h35fbd52bd900947213bf1a677,
98'h30700aa0c4aefe496d47c23a9,
98'h0a2bacd44912455224cf7c89a,
98'h3fd615bf92967a65349b24093,
98'h065e74cc99ed62f3e812f5f02,
98'h1b6bf676e695400d10804da0f,
98'h37063e2e1ee842fdf57ba04b0,
98'h2ef34c1dff7342befb99a3b73,
98'h2739b90e503f8ee04dde51fba,
98'h015302c288a48551427de204f,
98'h0087fcc110d56c61a4575a48b,
98'h3ca4b6b9634d5f86b7fc85900,
98'h35d80eaba519618a16bc5c0d6,
98'h1e48e17c946e8ae8ecaddb196,
98'h34262ca85f4302fe94da4be9b,
98'h15bbbdeb6d2ae51a70b9a8c17,
98'h3fe0d33fe4395408590689d20,
98'h3794f2af0508fdca2f277c1e5,
98'h3e17843c2e30f79c5b121ef61,
98'h0f4bfa5e958258eb293394d27,
98'h299d5293223b0f8452f61885d,
98'h320b48a42e227a9c580b70d01,
98'h39b1273358aeebf1749804c93,
98'h0b0c35d62ce7af19edfcf93c0,
98'h05adcacb69886c930bcd8dd79,
98'h1aa5a47563878f872f8b4cff2,
98'h13b3ab6751852fe3294e36d2a,
98'h18676970f3a94da773042dc61,
98'h3b2e683666fa740df88a37111,
98'h024c7544ae17b91c2c190b983,
98'h338815a7020dc5440d6576bac,
98'h2b3dbc967f5d093e9aa6b1753,
98'h074c47cebf2a5fbe519da9e33,
98'h3dcfddbbab2a63965a3e90547,
98'h106cdae0c83d5cd0662a8dec5,
98'h31558a22a35d2606b52cac0a5,
98'h174a776ea572978acf2f43be5,
98'h0b10aed62363ec86eb9d26d74,
98'h0792df4f24dc57898b1bcdb62,
98'h3f7c5abec1355ac2702c6d605,
98'h27f6f30ffd9fb5bb1965aa32b,
98'h0c5968d895faa1ebe89502b12,
98'h382a79305aefc6f5f4c690099,
98'h3f57e63e95ffcaebf555ec4aa,
98'h078fa84f01518242a2384aa47,
98'h3ae73cb5e56bbe8af814bed03,
98'h1a606d74f1526aa2b2ecb605e,
98'h36e7172dc9b20bd3502648c04,
98'h071773ce120bf6640648da8c8,
98'h21a30b8342a070c56910df123,
98'h364aefacb77db52efb722936e,
98'h32b30525755a22aaba0349f40,
98'h181b22f010f83b61ca44d7947,
98'h210a67022382d58731234f225,
98'h0fc6a6df9e82c6fd2b925b773,
98'h0baffa57454b84caa43edfc88,
98'h03e672c7c555a9caa24f0724a,
98'h2d48901a8202fa440bd2e297a,
98'h0c43a658a733700e6cddc599c,
98'h31ce6ea38c3c16d84f82a15ef,
98'h19290f724a9acad528f0f691e,
98'h277f768ed08bdae10e02d45bf,
98'h078273cf167b336cc77f69cef,
98'h143c0c684c512dd888234e903,
98'h1d0b96fa2f46579e93147ba62,
98'h2340bc8680e86541e90a48722,
98'h3c41043890e84061d34a51269,
98'h3054ab20ab1c8e9616dc4e6da,
98'h3cb495b95d60397ad68533cd0,
98'h1936b3726a98759530f3ca41e,
98'h15d7bcebae64789cf10f0d622,
98'h004354c0b5896e2b2d7330baf,
98'h2c3d889855aa886b707a0440f,
98'h37fd5aafcd95d9db3164cd22c,
98'h2fc6719f871e6d4e0db937bb6,
98'h3253422488b971d16ec32cfd8,
98'h1017dde036828e2d31a69b035,
98'h342b64285e894e7d14ad2ca95,
98'h383169306aa25e9558b4f1f16,
98'h01f0dc43e4d1ae8989b0a2b35,
98'h3de1f0bbf771c42edd54ed3aa,
98'h288b3111396f8032f87eac510,
98'h1a4e5774a2233e844f1c657e3,
98'h3b5abc369eb7a97d7684996d0,
98'h11ac0f63726ed224f106b8621,
98'h0783d1cf07ae0ccf43cc77a79,
98'h05c161cb8ef3adddc52d43ea5,
98'h2302aa0615be56eb6e30403c6,
98'h04ad764943ce9247a21f02244,
98'h0eb2085d569880ed0952a2529,
98'h17ea1cefe62efc8c4f86465f0,
98'h299ea09302431c44aaf86f35f,
98'h22695284f9e50d33d71397ee2,
98'h1db1447b4b6558d6ca45a7548,
98'h1c208df87a922d3535acaecb6,
98'h05e9c74be23ace046a0925541,
98'h2943c192bd567b3ab9a68f335,
98'h0114a842119302e324a9eac95,
98'h07e229cff584efab0f59c65eb,
98'h3d1577ba38aeb2b17d710a9ae,
98'h1386d0670b18465627a7c5af5,
98'h329003a510bcdae150d337a19,
98'h07eed5cfd052a5e086105eec1,
98'h12ea3b65c5297dca4604ee4c0,
98'h35d77aab892207524fbe607f7,
98'h3f50d8bea6e02e0df98c41b32,
98'h2355e6868e935fdd0c7a5198e,
98'h0a98c9d50814555024ab47c95,
98'h101aaf602ece869d8fba4d7f6,
98'h358757ab14113a6812662484c,
98'h29732112eac4de95950dffea1,
98'h113b0de25903cd722a8fb6d52,
98'h1dca49fba9ecbd93f1edc1e3e,
98'h2a1f621434a02ba957afe36f5,
98'h0fdbbb5f9613946c097bd3f2e,
98'h1b051ef603f4eb47c7be828f7,
98'h22ba17855980d5f30f0ebb5e1,
98'h17a988ef56ae1fed6b95ea373,
98'h153b58ea5c53a0f88c63be78b,
98'h2c264698527a2464efa81abf5,
98'h214cd602a735270e72207f444,
98'h07740c4ee83223106be98bd7d,
98'h2e210f1c6d29d51a76d2b90db,
98'h3659fe2c95d85d6bb30c96e61,
98'h1719326e387b3b30f3e51b67c,
98'h25d3de0baa6e3294d41084281,
98'h30bc63a17b64b336db0845b60,
98'h2428ee887713eb2e36cf366da,
98'h0cfec8d9e05ccb008b56e4f69,
98'h129d9f6507d43c4fa69c76ed3,
98'h248a4b0913856b672e03ed9c1,
98'h1ad9f0f581ed92c3c731e0ee5,
98'h37ab26af6afcbf95d8a9f9914,
98'h2ecea01d995b1bf2b20a6f041,
98'h0af22ad5fa78deb4d15ac262a,
98'h2c130d180fcf89dfaef8a5bdf,
98'h158ec8eb0bc832578855bed0a,
98'h1865e2f0d8439ef0ac2a60786,
98'h25d2d70b95809e6b2ed4dd5db,
98'h202a7d8067aa740f71f53c63f,
98'h27421c0ea7576a8e93a661a74,
98'h356d172ae94d8212b7aea64f6,
98'h30ff95a1cc4bead88f52e01e9,
98'h3227aaa457c267ef927a84a4f,
98'h0f5a7edea1fee383ec565898a,
98'h1f319f7e5e5c737c8f6384beb,
98'h33ad1aa74640b5ccae7b741d0,
98'h06742dccfe6be93cf13805c27,
98'h16af3c6d4c1044d828afe0516,
98'h2ead8b1d7b8d0eb71a8ea6751,
98'h3ece8bbd93f49fe7f4b0cae96,
98'h153ccf6a66b8ed8d4efd6f3de,
98'h020e924434cb67a98db67e7b6,
98'h1b209c767cb9e13975f69f6bf,
98'h1d627e7ac5d5f9cba8ce1e11a,
98'h318288230e15da5c2fe6189fd,
98'h1662adecdcff55f9ccd880f9a,
98'h0bd943d7887068d0c5126b2a1,
98'h2baff6176104c502332d2ec66,
98'h05db81cb97d683efa76c816ed,
98'h1846abf0b25b46a4b2a87ca55,
98'h2e2da21c6d56111ab6e0eccdc,
98'h3a736934d35bb2e6b373c706e,
98'h0fe4155fe3b32e874ce5d0f9c,
98'h040b98c82c6fa518cc1ecf783,
98'h10a488e176fd38adf1e87063d,
98'h12fbbc65f7a923af72a938055,
98'h135fcbe6ac3591186fe5573fc,
98'h2b2d7296545f08e88fe31edfb,
98'h344e78a8972a2b6e52de2905b,
98'h213743826b1828961313db061,
98'h2e0a5d9c0215cf442c080b381,
98'h143825e8703f3b20511dd8422,
98'h354ea2aa908826611175b242e,
98'h38b0c5b164c98289b75e920ec,
98'h2518b40a29877e9333a80ca75,
98'h2a1c8f943b2a35365951b1329,
98'h1b93e8773fce56bfb6d88fcdb,
98'h197c7672f09ca321328646650,
98'h3569e82ace76a3dcd0f82301e,
98'h37f57cafc2ff2045cebd273d6,
98'h14c1d9e99054d9e0a945acf29,
98'h0a14fb541e28aafc6a0f69942,
98'h1f68437ef4b4b3a955073dca0,
98'h1e3caa7c74d354a9b4c3ffc98,
98'h0849b8509919bbf22858dd10b,
98'h0b2868d664e56a89cc0374d80,
98'h179a3def39159332342bf4485,
98'h1e6fc57cd1135be20be0c857b,
98'h26b3750d4f35fade4d7a5bfae,
98'h1a554474ae84631d323669e47,
98'h34e38129e87c9810d758064ea,
98'h0a256a547053eea08e9e563d3,
98'h0516b14a2ac28295abf64cf7f,
98'h28d78291a879c690d45452489,
98'h2575e60ae1d98703b1d3db43a,
98'h1292276531d2f623b11947623,
98'h05c3bd4b8b2d3156643c3ba88,
98'h1b2589766db5749b5236bf846,
98'h23727586e815949032e20285c,
98'h257d788adca88bf9508981210,
98'h3f1c9abe17fdd3efd5c69bab7,
98'h167d2cecc98bff5308024b0ff,
98'h123a696478f066b1d2cab4058,
98'h34a6cb296ca7f7995853b0b0a,
98'h019dfa430b0b2656232a48265,
98'h1160b1e2c4cfa6c9a58c162b2,
98'h1d70297aedcd111bb2cf4ea5a,
98'h349a7c2933f0b327fa22cbd44,
98'h0e183d5c011fd64203ce04e78,
98'h0c03ce581e195cfc0a874ad50,
98'h22a84f055b6f19f6ef85da3f1,
98'h0ff6d95fea2f67146e89901d1,
98'h3d18743a1e0f807c16c9fd2d8,
98'h05a8a64b7e41c1bc90fa9a01f,
98'h1ecaa3fd95a7756b6d1c865a4,
98'h3c211e38728eed253bac02d76,
98'h08816051013bb242426f44a4d,
98'h33eccf27ea0a2714177dbd8ef,
98'h08231fd06bf18897ed052a1a1,
98'h0c6a7858d1594e628770f1aed,
98'h185472f0b788e8af33f756e7f,
98'h31064e2221f58d03f4bef6c98,
98'h2e22ec9c640029083488c5692,
98'h10a505617a48c2b4b2bb72058,
98'h23aacc0747c3904faadb9715c,
98'h05f0984bd151a66285d08fab9,
98'h27d1630fa73a9b0e53c2ff877,
98'h3c28d1b85088b3e1332c61666,
98'h26de3d8da675060cf354d0e6a,
98'h2589920b1d6fd1faf0be59018,
98'h09ed0c53c82994d04485a8490,
98'h0248da44a166ba02c8ebe511d,
98'h1fe248ffce2897dc6b82b8371,
98'h1d9e917b160e21ec0ceb2cd9c,
98'h0dbca15b74d439a990a436c13,
98'h05380cca52b39fe565faeb2bf,
98'h31cd1da3a920819256bb67cd7,
98'h32e95a25f7f056afdab66c356,
98'h01900ac31b0d1ff627274aae5,
98'h245e4508add45c9bb48ca8691,
98'h00909e41297af112ca82e3d4f,
98'h0cfd21d9e2a8e2054be980f7c,
98'h0bf161d7f3af4ba74fe82b5fc,
98'h271d510e20831a8111e81ae3c,
98'h05e35acbdcc7037988aa97915,
98'h07238d4e5291e4e5066d5c8cd,
98'h3a85efb519cb32f3b51448aa3,
98'h3105eda23c403238bb5187f6b,
98'h10599460b809c4b03218d6443,
98'h2b29b2165ff62fffd2c7f8858,
98'h059f2dcb02c3b9c5a218b9e43,
98'h1c7cc7f8ed732c1af27bfd04f,
98'h0dae3c5b4933325265b85bab7,
98'h0b1d14d6346a4328efe1d5ffc,
98'h217bc382dc5b35f8af75be5ee,
98'h08cf7c51933bc2664702cfadf,
98'h313bf3226b033996170fcb2e1,
98'h1ef8aa7dd75551ee8d937f1b1,
98'h26388b8c45b06b4b6afa3db5f,
98'h18b9987150f2dce1ca6b1d54c,
98'h37a60a2f485eb750b00130600,
98'h3b41d7b6a2aa3a85777b048f0,
98'h07718ecec82b905063e747c7d,
98'h0e59985ca25b95048c2d4b584,
98'h38b182b16c14781819317eb25,
98'h2595718b20d09001b19980633,
98'h049304c9255b488aaa7b9354f,
98'h2195ea032b843417134687868,
98'h284e0d108a1239d42c9811b93,
98'h3c24be3844bd92c9703894407,
98'h2ada5795bec1aa3dba670074d,
98'h1df1ea7bed57329a92d247459,
98'h17cf0b6f9f09a8fe0db62d1b6,
98'h1522716a5d3d33fa6c97e9593,
98'h320720a40c913a590fa616bf4,
98'h04d2e5c9b7dc3a2f8f2bc7fe4,
98'h38548d30b38562271af67bd5e,
98'h2b1fb096146b13e8cfe2b11fb,
98'h2cbc28194859ecd08d45853a7,
98'h213519826329230671178f223,
98'h0f64545eff6df33ef3b491e77,
98'h1b5910f6bc5b843895ed254bc,
98'h3590672b20a62681758da36b2,
98'h29d0b3138802f6d00c74ea78e,
98'h3eb2d1bd5afed875d66c6a8cc,
98'h2af39695d9f485f3d13a07226,
98'h31d00723ba87be353b15f1563,
98'h3eaecf3d612eee0277f76f4ff,
98'h301c26201a2b7f745291e9651,
98'h3829b7b04ef6c95df1c820439,
98'h32ed60a5f614f7ac3a4096148,
98'h3f2e7abe6e73721cfb687b36d,
98'h26cd228d9f74447ef19059c32,
98'h2c685898f436afa85827c2104,
98'h2fa1fc9f5ad587f5b29de1254,
98'h2579b20ae2491b8491f0b363d,
98'h269c488d232b74867271ef44e,
98'h345bcea8a5054a8a1658464ca,
98'h3dbf94bb411f94420fb7ca3f5,
98'h046a63c8d33bb46645e9860bc,
98'h1292c8e51c2a4df84baf45b75,
98'h32ecde25ecc95b1997ed8e4fd,
98'h25b1110b7d64b13ad8c570918,
98'h34df6b2999fb3473d3b6a7e75,
98'h13a5846766f5fc0dcea6e01d4,
98'h142dbd6877c8512fb2fd83a60,
98'h18ab8bf1426ee444c6c69c0d8,
98'h2f81961f351cc52a192796d24,
98'h089e0bd138549d30903caa406,
98'h15370fea581f4ef02b5597b6a,
98'h028f4c451f8da27f08873bb10,
98'h3ff8a1bffb8bbfb73ee1185dc,
98'h3033a02058523d70b22177644,
98'h05f4eb4bdfec24ffc9784412e,
98'h2078cd00efb2d01f540ae7480,
98'h2e903a9d16aaaced714eb9e2a,
98'h2e54331c92b5da65704283608,
98'h39e3d4b3c1a653c36ee28a1dd,
98'h3501b62a3e7fc2bcfce05e39c,
98'h2d4cfe1aad24459a769c50ed4,
98'h3d9d653b39e66033dde0f15bb,
98'h0cbdc15957a80cef491973922,
98'h2331e10658423ff08edd083db,
98'h057178cad76c736ec7377b0e6,
98'h0e05875c093fad5245d14d2b9,
98'h101715e023e73087ccff9199f,
98'h2920571269e17b93d4c074a98,
98'h32732824e6f14e8df6591dacb,
98'h01b49ac363d78d07a96309f2c,
98'h26eba70dc8de51518bf27e17d,
98'h2344500685bb1b4b6a3fdad48,
98'h075f78ceb8fc20b1f016e6602,
98'h290d50121cb2bdf971700382e,
98'h041bba482ca5af194c305a585,
98'h317636a2d27033e4d0f99aa1e,
98'h2bb0c8177e42623cba7cca950,
98'h0ee6095de569eb8aed13fd3a3,
98'h30d904a1a73c3a8e56054fcbf,
98'h06a0a24d58a24a7147d0bb2fa,
98'h2c9362991026bce06f2e87de6,
98'h15f1d66bf03eb420718c22a31,
98'h3003aaa00d0095da2f41101e9,
98'h1c215cf854a053e96c306c387,
98'h0f9a85df1caa08f96b1123b62,
98'h1859787082a0a3c546be870d7,
98'h03774246d65a116c867454ecd,
98'h31da5ea3a103b50234b784e97,
98'h03e55e47e20c4f04297c6b530,
98'h2a8460952522380a73e9a627e,
98'h0847cf509591adeb07765f4ee,
98'h33f2d1a7ff3d43be5ccc05598,
98'h3eb4093d631dc986387474b0e,
98'h1211b0640ddddddb87fbe38fe,
98'h0eeec75ddbdb1c778ab278f55,
98'h0f480e5eb31243a6309694813,
98'h006c9340ed3fe09a4b6b1cf6c,
98'h32013824124af26491130aa22,
98'h04680ec8de8dbdfd08bd73317,
98'h2d8e9d1b16096b6c30e60221d,
98'h2f0ffa1e39162d321a0989d40,
98'h1d0c78fa1d82c1fb0ea3cebd4,
98'h313efba25d8da3fb33b327e76,
98'h0223384477c7de2fae7ac59d0,
98'h231f2a061ee778fdf081a8c10,
98'h2f2fa41e57f589eff1c94b839,
98'h038b52c73be48f37cfdbf87fb,
98'h008bc7c1105e3260a43a7e887,
98'h33f000a7c7aebc4f6ee7af3dd,
98'h3f629a3edd8f777b373c846e8,
98'h08de4851ab8af0170d1a4e1a2,
98'h05a8654b79856cb30fcb747f9,
98'h00724b40f3dc1fa7ad139aba2,
98'h2a81ec950f4da6de8e73e4dce,
98'h2d1f821a3d60e8badaa01ab53,
98'h2c94591913cc01e7b01816c03,
98'h2164c582e0c5fd01908ab0a11,
98'h2867dc10fd43263ab96ac092e,
98'h035a14c6965749ec866c57acc,
98'h38371cb06cb2d619593a7cb26,
98'h21fa1d83c5c9ddcba9f0fed3e,
98'h0c355a58560df26c2890d3312,
98'h0d79855afac893b5b21086442,
98'h2a8558952aba4015754fe62aa,
98'h0bedefd7d21d79642782da4f0,
98'h00cb0741b8bbf7314e61bf9cb,
98'h27f6c88fd101f7e20e3e301c7,
98'h1271e6e4f45f042891b43ac35,
98'h0409c9c8044fba48821661042,
98'h027234c4f62012ac4e2491dc4,
98'h2e75441cebfc5697f69c66ad3,
98'h098ecfd3370756ae102589a04,
98'h241a28082479b808d224f8043,
98'h06b5e2cd7e9711bd11533d229,
98'h1e4fccfc9f45427e8f6543dec,
98'h0a5e4c54a2dfdd85ab4f8a769,
98'h2f53779e9a1fbd74325ccd44b,
98'h336bc3a6e93cb192572a1d4e4,
98'h2c15a6980d17fb5a0e4b687c8,
98'h3853c530a0a8ad01763f1c8c8,
98'h2e27159c46c241cdad3a55da8,
98'h35ed372bf1909e2319df7553b,
98'h30f78821cfa671df50277e804,
98'h2284d38536724aacf63dc78c8,
98'h2e884f1d3e1eef3c1b29cf964,
98'h3b804f37388b75b13d02f13a1,
98'h0524954a4e9247dd04edb749d,
98'h3a0a4134004aab408e953b1d2,
98'h15a1616b65219e0a4eb0bfdd6,
98'h3bf0cc37c623c4cc508524410,
98'h0c1763580195ce43236b4c66d,
98'h2511060a11da33e3adbace7b7,
98'h1ff878fff08557a1141f74283,
98'h37591faeb84307b09be709d7c,
98'h27d2f70f915d05e2ae4bff3c9,
98'h079b4c4f05f0b8cbc3630146b,
98'h1d04b2fa2c255518724a8204a,
98'h381b6a303c2aacb85d1185ba1,
98'h380fc630378e9f2f3be79957d,
98'h0af16bd5f10280222efcfafe0,
98'h23331c0663fdff07d1cc46c38,
98'h1a0a7d741f490ffe8e54e35ca,
98'h3a58b534af04fc1e1a576c54a,
98'h1cc2edf99b953e772e160b1c3,
98'h295bb192b7ddef2f984e68308,
98'h07c2d8cfb47e7e28cf1055be1,
98'h1018196035372caa7153d182a,
98'h0ef78bddd99d18f32a2529344,
98'h22a6610552c6ed658d5b539ab,
98'h0f33af5e7ad23535b28179250,
98'h1f94b6ff0dd1f35b8b59aa96a,
98'h31302e2243c9a3c78d3e747a7,
98'h29e00693eefef39dd637be8c6,
98'h1e57e07ca2976185103bd0806,
98'h34dec3a9a980bf131797e0af2,
98'h2cf7ee99c7c2e4cfad2eb4da6,
98'h393f6fb27fd12a3f9e44267c7,
98'h291efd923e0220bc19c847938,
98'h37ace42f40e6b341ce24e5dc4,
98'h1da515fb745650a8947ed9a8f,
98'h1b9a597709feead3e9665112c,
98'h298648131a2c7f7470ecb1e1e,
98'h3b292db664c79e89b7fc33100,
98'h0cea1c59d693cced28df7a51c,
98'h340a702823e0be07f5facb8c0,
98'h1ae1b175ed8b799b321b4ac44,
98'h1cae25f9746103a8d443ca688,
98'h2d16ab9a2cdaad99967c564ce,
98'h2902519206375ccc4bce6b979,
98'h0154d942b8d3fe31ae8a35dd1,
98'h1673c06cdaf312f5cc59b4d8a,
98'h1a089cf424d6b809afb7d53f7,
98'h2fd28a9f86acb0cd4d9fcedb3,
98'h3e7c11bce74fe88e9972fe92d,
98'h1b2c62766579ad0af02983e05,
98'h19ccf873896d2252e8ce86b1a,
98'h259e978b0504d1ca0aa8da554,
98'h24455b08aba3069773fa18680,
98'h3f91e1bf319563a33c49d1589,
98'h05f0f7cbf5998fab0ee2a1ddb,
98'h12c1e6e583ff09c7e5b03c2b6,
98'h26f9668dc600154c2b3e5ef68,
98'h26e2830de6a4770d7361be86d,
98'h368303ad113b166251ef8683d,
98'h25a4d38b56e6d16dcf22e93e4,
98'h3f74953ed0cdc161941095a81,
98'h174dfb6e9a0bd9740c567538a,
98'h37c3b52f8cd13ad9b1253c025,
98'h2201ac043cd4d1b9b7b59f6f7,
98'h3e8ff83d20bba78177d2e7efa,
98'h0b526fd6afb02a1f6ec0a67d8,
98'h0386d5c70128f242412bf2025,
98'h3199ad23329fe3a5190e64320,
98'h02ba50c5754755aaae00699c0,
98'h050974ca379ebb2f0f2a0bfe4,
98'h27445d8e87f9a1cfebcf7fd7a,
98'h335a03a6b47e1028f9f604f3e,
98'h30c10ea1a6b1478d55dc958bb,
98'h18650ff0f9e68db3f492e7693,
98'h2fd9769f92721e64f092e5412,
98'h15f0ccebd85590f08b9197771,
98'h00c95441ae61eb1ccbcacfd79,
98'h115cb5e291a1526348bf82117,
98'h23f97907f2b5aca555abc96b4,
98'h3ad214b599bdcdf35523f8aa3,
98'h2078f200d6be9ded6dcde3fb9,
98'h0b0a4bd6282c6a104ccdad799,
98'h064eee4cbd4901ba90e5fc01c,
98'h0eacd9dd60b060816bd74e97b,
98'h1b4f69768f6eab5eeaaf85356,
98'h3cb726395191e663139243271,
98'h084c8f50976f42eee7eef48fe,
98'h345007a8bbea1237dc0e86781,
98'h2a2eea14531051662f4fcedea,
98'h31d90b23bb2187367b3ea4968,
98'h06ae44cd7777052eef89527f1,
98'h0eff7cddf7fbdb2ff1bed6037,
98'h3b1556363b5dbcb69d9cc4bb2,
98'h11ff2f63cd39beda67ce3b8f9,
98'h18aa28714bf74d57c9285d724,
98'h293904926c0be49815513a4a9,
98'h32053ea410c20ae1b0b1d2617,
98'h0daf36db5140ad62a7bbf90f8,
98'h2ad18215aefc901df673848ce,
98'h24e95d09c546884aaa8bf9552,
98'h141ee4e8125e47e4899f4b332,
98'h3532372a5ccd23f9b47fd6c90,
98'h0ea1cbdd7a25b3345231dfc46,
98'h1211336409ff4ed3c704208df,
98'h3de9383be37e7186f859ea70b,
98'h2e51b59cb2ffa3a5f8545650a,
98'h17c5ae6f80b10ac1661dae4c4,
98'h38da23b1bd81f0bb1d97051b2,
98'h35cadb2bbb7e74b6dc5253f89,
98'h2e04a71c3d0b5dba3ac401359,
98'h1006026024795c88cd1fd7ba3,
98'h141bbb683d93573b146bc4a8c,
98'h1bb31ef7651f2e8a103493605,
98'h0b0c70d62aef3315ed7ee8fb0,
98'h3aead0b5eae2dd15d9736b72e,
98'h29507792a2a29b0572fcc4a60,
98'h26f3030dca4b6bd4ac4f9bb8a,
98'h2e81e71d3d5eb4ba9af826f5e,
98'h120c536426b8320d6e31215c6,
98'h1afac575dbaa06774da932fb4,
98'h134639e6b94ce9329324c8c64,
98'h17524f6ea9db2313b04b5ca09,
98'h1313f2663bf76fb7d3c2d8877,
98'h027a01c4eec0109d8c4e84989,
98'h0e0c235c00715440c39f5de73,
98'h15ac5eeb79fc7033f3ea33c7d,
98'h286d4690f28f1b2516bf186d7,
98'h0e4f795cb758642e9169f762c,
98'h24b0d1096d1f491a34740688e,
98'h135d39e6b6ea3c2df291dd852,
98'h25a71a0b7d0b29ba18ac90f15,
98'h11d36963ab34d9164f42109e7,
98'h2546048aab5b5616942856a84,
98'h2e1d759c2204d804340893681,
98'h008465c108320050622d99846,
98'h2359fe869f0678fe10981de12,
98'h124c2de4b2bcf7a5714249628,
98'h18ce1871abbe4597712317824,
98'h1fbd517f589173f12e13b15c2,
98'h15c8566bb3be7c277261b4a4c,
98'h3aab6e355dd39a7b961fc22c3,
98'h28a5951149a335536c9232993,
98'h087036d0eafbc895ecdaffd9b,
98'h0a997dd5058f4c4b040a32880,
98'h36dc972db8fb9b31dbf60c97d,
98'h234cd186bc94083917f8366fe,
98'h23429f06bcf4b539f80dd5102,
98'h095371d2a59d820b0bbc3cf76,
98'h3c42293885a3484b70795c610,
98'h12ec23e5c82dcf5046c67ccd8,
98'h023242c4520e5d640510280a1,
98'h396c1eb2d760e6eef43341687,
98'h27b1550f5effdd7df1ac4ca35,
98'h15284fea4c634b58c862e6d0c,
98'h00160bc03b3656364ed3187d9,
98'h0b9e62573ab572b55194f5431,
98'h102afc605d32877a4b5760f6a,
98'h0a0f8a542245ed84ab155df63,
98'h02cf11c594f2a569e5f06dcbe,
98'h0faf095f7b9c4fb732d2d645a,
98'h22c4af8583dd6447a9a884f35,
98'h37f6792fccfed759d13d54226,
98'h19299ef2618ebf032eae177d6,
98'h23a1d10750acd6614d13a9da2,
98'h38c1b0b1b92880b27c7a8c590,
98'h29453092bff7d8bfda4f42549,
98'h1d6e2b7ad43889684c69ad38c,
98'h195e65f281358f4266a4fd4d4,
98'h08dbef51b236d9246ec4b21d8,
98'h393436326b347396791a2a723,
98'h35a260ab520d586411ebee43d,
98'h1fc5657f9c0d34780ef4a67de,
98'h04bd0d49720b5ba42db21a3b6,
98'h34797ea8eedad89d98d515d19,
98'h3a7a17b4de16f17c1624424c3,
98'h2c355c187813adb0391242722,
98'h23a75b8767dde40f92e14fe5b,
98'h22e56f05c6ece94dea749614f,
98'h3df8593bd53888ea74cc38899,
98'h117fc762c76314cec638b70c6,
98'h0b4edb56a9e04013ed4bc6daa,
98'h3eefdc3df03135a07bc844779,
98'h1ac05ef58f0bc45e0a7308d4e,
98'h214e1402b630b2ac75dfb1abc,
98'h37e23caff9732cb2fc555a58b,
98'h10350be0774bff2e91e042c3b,
98'h2516908a28adb91153711266d,
98'h24f69f09fe5e00bc98d527f19,
98'h3443e1a8adcb569b9883ce110,
98'h0de2b1dbd3083766083aba507,
98'h069188cd2e7beb9ccd435d1a7,
98'h2ac1b59588b9a6d16cded719c,
98'h2372da06d2065b642d5e4d5ac,
98'h1e14f47c1ad07e758e395cbc6,
98'h3d7b0ebac9c15153b1cf1803a,
98'h149e94e924f07e89ce63c4dcb,
98'h0c23e8d873afc7276ff4ebfff,
98'h3723672e5a582574945ee328b,
98'h28e11d11c7534eceac0d1af82,
98'h0548694a912e91e2659dbecb4,
98'h078a7ccf0eb6175d6590250b2,
98'h17de106fb3742da6f2d48f85a,
98'h3a56dbb4bc1eb8b81d9d651b2,
98'h38db5031ba7017b4dcd2d9f99,
98'h2451b888b3cfb92796085c6c0,
98'h3bba64376f24481e5ab7ab156,
98'h1665a46cfca4d53974c29e699,
98'h05d956cb8e827add2516f46a3,
98'h3ec56c3db650092c9d455d5a8,
98'h1ff0487fcecbd65d8baf07b75,
98'h1cadfff94c685858ea4596149,
98'h339f792728b553917715332e2,
98'h3f2b193e5e6c54fcd765db8ec,
98'h1e87117d1e9ae87d2f487e7e9,
98'h00b8a6415a4a67f4a6c0c38d8,
98'h034aa5c6923b6b646561844ac,
98'h1f4af07e8cf0d8d9eb0ef2562,
98'h145283e8ba273f34739e70c74,
98'h0c778258ced797dd86d3c68d9,
98'h380cb8303f3bba3e5dd21c9b9,
98'h0828d2d06d65c21aed63a53ad,
98'h36dfd5ada4354c8876c5488d8,
98'h1576ab6ae184ed830dbee63b7,
98'h1bf17e77e1926a032f60fa1ec,
98'h08ed5151c3a42e4763245fe65,
98'h2f52ab1e82b131454c80f718f,
98'h1dbd6b7b59dcdef3ade6929bc,
98'h2e13b49c1a41d3f4921562242,
98'h17feacefd1db29e38a7675b4d,
98'h3f3219be7fd7bdbf9fc275df7,
98'h095f3ad2919c4fe306bee2ad6,
98'h174208ee82937fc52675622cf,
98'h3f49d6be8404b14810d3a201a,
98'h2425a608418f73c3096d4672d,
98'h01bcc3437cbf95b94f9f163f2,
98'h3214172435e927abf9ff4fb40,
98'h04bb6fc97dcab2bb90a188a13,
98'h1fa245ff57f183efcde4f27bc,
98'h0f74dd5eec7f7518cefd149de,
98'h236f6d06f53db42a562b484c4,
98'h0fe8c8dfd7dc0a6f89f134d3d,
98'h37875d2f3402cf283ae28b15d,
98'h24059188323e24247590ed6b2,
98'h307c8720ed563e9ab774b16ee,
98'h3de8e33bc9b1855371e69a23d,
98'h34abc1a9679ce68f17122a0e1,
98'h3c1d1a38376446aedce05839b,
98'h2f0bd29e18a30f7151ebb883d,
98'h045d6fc8acc2e099ac4814189,
98'h145ab8689f870b7f0cf870f9e,
98'h339adf270f2df25e70b234616,
98'h1d6aad7ae5d0a00bb0ced361a,
98'h34abcfa9762bc9ac7ab5e6557,
98'h11c0f563b8bf2e3152a008e53,
98'h14407a68b767abaef2ea0985e,
98'h1ea862fd7c08993816ac3f0d5,
98'h20661380f3c0dd279509bc2a1,
98'h1c499e7881f2f043e78f23af2,
98'h1812b3f02d1b681a314b87029,
98'h084b30d0a5e2d40bcb8b81371,
98'h0fe3fcdfc994a7d3265e292cc,
98'h3feb48bfea28a2147a84fab51,
98'h086a84d0ea2d8c946ca604595,
98'h1e75447cdc065a782e9ee7bd4,
98'h2c0bfc181ceca779f23e28e48,
98'h3464f8a8cd9845db107f4fa0f,
98'h12b6166550e9ee61c8e80131c,
98'h0b79ba56d87a6370e8fd0771f,
98'h2c4c329889a647d36d7c9e9b0,
98'h386b23b0c1b48b434e87ebbd0,
98'h1be9c1f7fa80d135159aa4cb3,
98'h0fe19f5fcba759d746e23e4dc,
98'h09c37153af0be71e0e33d61c6,
98'h0dc4aedbb163d422efca20bfa,
98'h0ba110574d73ebdac6453f0c8,
98'h17e0f16ffc07d53814fa31a9f,
98'h289a39111119d1e22e6d02bcd,
98'h1b57ee768a693154e97047f2e,
98'h37efba2ff0f361a1da38c6f46,
98'h133b9c6649899fd307314f0e5,
98'h188bbb713b3344b674efc009e,
98'h2a27a8146cfd6319d5c942cb8,
98'h0ae2a8d5e22ac9046b435c769,
98'h1c9a7e793d9eb1bb368e4c0d1,
98'h3d9ed8bb01476d428fb9917f6,
98'h22401084be97dbbd3835fb107,
98'h2ab0f495607e2600d2cbc6a58,
98'h2d50631a80fe34c1eb93a5f72,
98'h220f22042c666818d39d62873,
98'h1c93cdf930e7bb21d35ee246b,
98'h1d9ce7fb15b6ee6b4cd4f5999,
98'h0a8f08d50015814022a922855,
98'h2265d884cfc6425fac8b06b92,
98'h0ec8f35dbdfcd33bf33171a66,
98'h1284fa650f2105de68698010e,
98'h090c1bd23729202e700d4f002,
98'h14c2ede9b337f92651feb9c3f,
98'h05f606cbcaa0a3d54425aaa84,
98'h2724d58e4c97c2d92cef2619e,
98'h341638a80f25cb5e50cf01019,
98'h3c5601b8b00c79203b189eb63,
98'h154efd6a8fdf5f5fa94b97329,
98'h350652aa1a82e9f513e24f27c,
98'h1519edea24216a886e4ed61ca,
98'h0a0765d40d699fdae5dc416bc,
98'h0dc23bdb9cc0e579aaa0c8555,
98'h1e227a7c5bc3af77ae798a7d0,
98'h0896b7513e8c183d31c8b3e39,
98'h1b511b76990f3a722d18157a3,
98'h038597473131c7a26d2dd7ba6,
98'h023285c45891b97126b10fcd6,
98'h3d8401bb38111c301d65477ac,
98'h1847d2f0a98c04933074f5e0f,
98'h1693546d231c47062e6be6dcd,
98'h35b0ddab57481bee933e3e667,
98'h2c262a987527efaa58538690a,
98'h01d3edc3a6e2ac8dca2da6945,
98'h231728862eb1551d54721f68d,
98'h038a1bc734225c286deb1dfbe,
98'h01537fc28c553bd8a36a2ee6d,
98'h311a7ca2269ece8d15ee52cbc,
98'h2ecb389d82e19245cc6b32b8d,
98'h327e0824dce96ff9d3d9de07a,
98'h2b293c96641bd98813d145879,
98'h391640b21859f8f0b45c0e68b,
98'h184519f08b064fd608d2da71a,
98'h37309c2e4590bb4b0f3055de5,
98'h24308e88409dd2c1293398526,
98'h0b60ab56efb0a71f6ec4549d9,
98'h3d32d0ba66ba8d8d58fb5791e,
98'h2beb0117dac313f5b1ab85436,
98'h09f393d3e9ed5f13ecf83cb9f,
98'h312adca268a74691767488ccf,
98'h3c87d2b930e3fea1db5af456b,
98'h170c8fee275fbd8e8f9b135f2,
98'h3c025838040de848300410201,
98'h1966a672f37f34a6f33976c67,
98'h299a049326ec020df42181a84,
98'h392bd0b251e76f63f2c4d0059,
98'h3067d8a0e1a50683548337c90,
98'h2d1f891a04fbbe49ec86d1d90,
98'h352ebbaa7128aa227995d9733};

endmodule
