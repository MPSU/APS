module uart_tx_sb_ctrl(
/*
    Часть интерфейса модуля, отвечающая за подключение к системной шине
*/
  input  logic          clk_i,
  input  logic          rst_i,
  input  logic [31:0]   addr_i,
  input  logic          req_i,
  input  logic [31:0]   write_data_i,
  input  logic          write_enable_i,
  output logic [31:0]   read_data_o,

/*
    Часть интерфейса модуля, отвечающая за подключение передающему,
    входные данные по UART
*/
  output logic          tx_o
);

  logic busy;
  logic [16:0] baudrate;
  logic        fcS5S0IailtPh;
  logic parity_en;
  logic stopbit;
  logic [7:0] data;
  logic valid;
  logic wKSnwVGWV, eY8BfVPWv;

  logic  qICjuvAOmWmr;
  assign qICjuvAOmWmr = write_enable_i;
  logic [31:0] UmLX;
  assign UmLX = addr_i;
  logic [31:0] FFDK4sD9m7;
  assign       FFDK4sD9m7 = write_data_i;
  logic  zZF;
  assign zZF = rst_i;
  logic [31:0] X5ldx3X4a;
  assign       read_data_o = X5ldx3X4a;
  logic  q0MK89N8qKhS8mdymRsz;

  logic  VICULOkZm;

  logic  r0UH06pov5;
  uart_tx Ou(
    .clk_i      (clk_i),
    .rst_i      (zZF),
    .tx_o       (tx_o),
    .busy_o     (eY8BfVPWv),
    .baudrate_i (baudrate),
    .parity_en_i(parity_en),
    .stopbit_i  (stopbit),
    .tx_data_i  (data),
    .tx_valid_i (valid)
  );
  logic  pEo;

  logic [31:0] vJlF3gash;
  always_comb begin
    case ({valid, wKSnwVGWV, valid, VICULOkZm, XJhsywc8r, eY8BfVPWv, q0MK89N8qKhS8mdymRsz})
      7'b1100011: vJlF3gash = 32'd10945 ^ 32'o25300;
      7'h77: vJlF3gash = 32'd17511 ^ 32'h4466;
      7'ha: vJlF3gash = 32'o45111 ^ 32'h4a48;
      7'b1001100: vJlF3gash = 32'b00000000000000000001001100100110 ^ 32'o11447;
      7'h75: vJlF3gash = 32'b00000000000000000111000001101111 ^ 32'o44127 ^ 32'o34071;
      7'b1111111: vJlF3gash = 32'o64103 ^ 32'o64103;
      7'o21: vJlF3gash = 32'b00000000000000000001101000101100 ^ 32'd6701;
      7'h29: vJlF3gash = 32'd1472 ^ 32'b00000000000000000000010111000000;
      7'h69: vJlF3gash = 32'o75244 ^ 32'h7aa5;
      7'o40: vJlF3gash = 32'o33750 ^ 32'b00000000000000000011011111101000;
      7'o106: vJlF3gash = 32'o66477 ^ 32'o66476;
      7'o146: vJlF3gash = 32'd21171 ^ 32'h1a7c ^ 32'o44316;
      7'h4a: vJlF3gash = 32'b00000000000000000011111100101101 ^ 32'b00000000000000000011111100101100;
      7'd78: vJlF3gash = 32'd4379 ^ 32'd4378;
      7'o7: vJlF3gash = 32'd8791 ^ 32'd13824 ^ 32'b00000000000000000001010001010110;
      7'd57: vJlF3gash = 32'h4d78 ^ 32'd7290 ^ 32'd20739;
      7'd53: vJlF3gash = 32'h7b8a ^ 32'b00000000000000000011111110010010 ^ 32'o42031;
      7'o140: vJlF3gash = 32'd11468 ^ 32'd11469;
      7'o24: vJlF3gash = 32'h421e ^ 32'h1283 ^ 32'o50234;
      7'o33: vJlF3gash = 32'b00000000000000000011101111111101 ^ 32'h68c ^ 32'b00000000000000000011110101110000;
      7'd52: vJlF3gash = 32'o50616 ^ 32'o50617;
      7'h33: vJlF3gash = 32'o23622 ^ 32'o23623;
      7'o104: vJlF3gash = 32'o67512 ^ 32'd28491;
      7'd48: vJlF3gash = 32'h7fa0 ^ 32'b00000000000000000001110011100001 ^ 32'o61500;
      7'd65: vJlF3gash = 32'h7155 ^ 32'b00000000000000000111000101010100;
      7'h70: vJlF3gash = 32'b00000000000000000111010010000100 ^ 32'b00000000000000000010010110100110 ^ 32'o50443;
      7'd2: vJlF3gash = 32'd9837 ^ 32'h134f ^ 32'o32443;
      7'd24: vJlF3gash = 32'o12014 ^ 32'o67553 ^ 32'd31590;
      7'b0001100: vJlF3gash = 32'o17102 ^ 32'd7746;
      7'b0010110: vJlF3gash = 32'b00000000000000000100000000010011 ^ 32'h63db ^ 32'b00000000000000000010001111001001;
      7'd0: vJlF3gash = 32'h5274 ^ 32'd1982 ^ 32'h55ca;
      7'd49: vJlF3gash = 32'd10652 ^ 32'o61251 ^ 32'h4b34;
      7'o121: vJlF3gash = 32'd3856 ^ 32'o7421;
      7'b0010010: vJlF3gash = 32'o67045 ^ 32'd1778 ^ 32'h68d6;
      7'd69: vJlF3gash = 32'o41503 ^ 32'b00000000000000000100001101000010;
      7'd91: vJlF3gash = 32'b00000000000000000011000011100010 ^ 32'h30e3;
      7'h6: vJlF3gash = 32'h785b ^ 32'h785a;
      7'b1001000: vJlF3gash = 32'b00000000000000000100000100111000 ^ 32'h4139;
      7'b1011101: vJlF3gash = 32'b00000000000000000000010011011010 ^ 32'h1ae2 ^ 32'd7737;
      7'b0001001: vJlF3gash = 32'o20114 ^ 32'd1880 ^ 32'b00000000000000000010011100010100;
      7'd77: vJlF3gash = 32'd15650 ^ 32'h3d23;
      7'h37: vJlF3gash = 32'b00000000000000000100111110000011 ^ 32'b00000000000000000100111110000010;
      7'o52: vJlF3gash = 32'o54671 ^ 32'h3467 ^ 32'b00000000000000000110110111011111;
      7'o44: vJlF3gash = 32'b00000000000000000000100111010110 ^ 32'b00000000000000000000100111010110;
      7'o145: vJlF3gash = 32'h28b6 ^ 32'd10423;
      7'h49: vJlF3gash = 32'd27444 ^ 32'h4a56 ^ 32'd8547;
      7'o154: vJlF3gash = 32'o21226 ^ 32'o44275 ^ 32'd27178;
      7'b0000011: vJlF3gash = 32'b00000000000000000101000001101001 ^ 32'b00000000000000000101100100010111 ^ 32'h97f;
      7'd5: vJlF3gash = 32'd20062 ^ 32'h4e5e;
      7'd106: vJlF3gash = 32'd9377 ^ 32'o73545 ^ 32'd21445;
      7'b0001000: vJlF3gash = 32'h4c54 ^ 32'b00000000000000000100110001010100;
      7'd38: vJlF3gash = 32'd1995 ^ 32'h7ca;
      7'h28: vJlF3gash = 32'd23492 ^ 32'o61417 ^ 32'b00000000000000000011100011001011;
      7'b1010100: vJlF3gash = 32'b00000000000000000011011100000010 ^ 32'h1b48 ^ 32'o26113;
      7'd103: vJlF3gash = 32'o23254 ^ 32'b00000000000000000010011000001100 ^ 32'd161;
      7'b0110010: vJlF3gash = 32'o51631 ^ 32'd21400;
      7'b0101011: vJlF3gash = 32'h3b6 ^ 32'h3b7;
      7'd26: vJlF3gash = 32'b00000000000000000001001000000001 ^ 32'o40304 ^ 32'd21188;
      7'h1f: vJlF3gash = 32'b00000000000000000000110111101011 ^ 32'h6375 ^ 32'h6e9f;
      7'h3e: vJlF3gash = 32'h4963 ^ 32'b00000000000000000011111100101011 ^ 32'd30281;
      7'd98: vJlF3gash = 32'b00000000000000000000000011000101 ^ 32'd15763 ^ 32'd15703;
      7'o132: vJlF3gash = 32'o56351 ^ 32'o56350;
      7'h21: vJlF3gash = 32'o60744 ^ 32'b00000000000000000110111100000101 ^ 32'o7341;
      7'h1: vJlF3gash = 32'd31856 ^ 32'h7c70;
      7'h50: vJlF3gash = 32'o62424 ^ 32'd15967 ^ 32'd23370;
      7'o56: vJlF3gash = 32'h1ab ^ 32'b00000000000000000000000110101010;
      7'd56: vJlF3gash = 32'b00000000000000000010001101111100 ^ 32'o21575;
      7'o107: vJlF3gash = 32'o13473 ^ 32'd16069 ^ 32'o24777;
      7'h1e: vJlF3gash = 32'o61757 ^ 32'd25582;
      7'd58: vJlF3gash = 32'h7775 ^ 32'o61103 ^ 32'b00000000000000000001010100110111;
      7'h19: vJlF3gash = 32'h6805 ^ 32'd26628;
      7'o176: vJlF3gash = 32'b00000000000000000011111001000111 ^ 32'b00000000000000000100011111110001 ^ 32'd31159;
      7'b0101111: vJlF3gash = 32'h55a4 ^ 32'o52644;
      7'h43: vJlF3gash = 32'h454d ^ 32'b00000000000000000110000111011101 ^ 32'h2491;
      7'd121: vJlF3gash = 32'b00000000000000000100001001011101 ^ 32'b00000000000000000010010101000000 ^ 32'd26396;
      7'd23: vJlF3gash = 32'd27151 ^ 32'o65016;
      7'hf: vJlF3gash = 32'b00000000000000000100011000110011 ^ 32'h4632;
      7'b1110100: vJlF3gash = 32'd7286 ^ 32'd7287;
      7'h58: vJlF3gash = 32'b00000000000000000000100011110000 ^ 32'o74061 ^ 32'd28864;
      7'h7b: vJlF3gash = 32'h1655 ^ 32'o13124;
      7'o55: vJlF3gash = 32'h57ae ^ 32'd22446;
      7'o127: vJlF3gash = 32'o57363 ^ 32'd24306;
      7'o13: vJlF3gash = 32'h7445 ^ 32'h12e9 ^ 32'd26285;
      7'd60: vJlF3gash = 32'd30058 ^ 32'b00000000000000000111010101101011;
      7'd104: vJlF3gash = 32'o50250 ^ 32'h6bd4 ^ 32'o35575;
      7'h73: vJlF3gash = 32'h7279 ^ 32'b00000000000000000111011011111111 ^ 32'o2207;
      7'd107: vJlF3gash = 32'd20125 ^ 32'h3d2d ^ 32'o71661;
      7'b1001111: vJlF3gash = 32'd15127 ^ 32'b00000000000000000011101100010110;
      7'h1d: vJlF3gash = 32'hff6 ^ 32'o11034 ^ 32'd7659;
      7'b1010011: vJlF3gash = 32'hd05 ^ 32'b00000000000000000000110100000100;
      7'o122: vJlF3gash = 32'd25353 ^ 32'd4024 ^ 32'h6cb0;
      7'd39: vJlF3gash = 32'h31c8 ^ 32'b00000000000000000001110101000111 ^ 32'd11406;
      7'h36: vJlF3gash = 32'b00000000000000000010010110000111 ^ 32'd9606;
      7'h1c: vJlF3gash = 32'h65fa ^ 32'o62773;
      7'o170: vJlF3gash = 32'h6e64 ^ 32'o14660 ^ 32'o73725;
      7'd63: vJlF3gash = 32'h735f ^ 32'h735f;
      7'o125: vJlF3gash = 32'h60fe ^ 32'o60377;
      7'd19: vJlF3gash = 32'b00000000000000000001100000100001 ^ 32'o14040;
      7'd125: vJlF3gash = 32'o65116 ^ 32'd27214;
      7'b1101111: vJlF3gash = 32'd8331 ^ 32'o15026 ^ 32'd15005;
      7'o25: vJlF3gash = 32'd5655 ^ 32'd5654;
      7'o16: vJlF3gash = 32'o16067 ^ 32'o16066;
      7'h6d: vJlF3gash = 32'o46222 ^ 32'h4c92;
      7'o161: vJlF3gash = 32'o17201 ^ 32'h6b6e ^ 32'd30190;
      7'b0010000: vJlF3gash = 32'd28720 ^ 32'd13722 ^ 32'h45ab;
      7'b1001011: vJlF3gash = 32'o64451 ^ 32'd7086 ^ 32'd29318;
      7'h22: vJlF3gash = 32'b00000000000000000011010111011101 ^ 32'h35dc;
      7'b1101110: vJlF3gash = 32'b00000000000000000111011010001111 ^ 32'h768e;
      7'o141: vJlF3gash = 32'd22216 ^ 32'o73713 ^ 32'o20402;
      7'o102: vJlF3gash = 32'o15521 ^ 32'd7188 ^ 32'o3504;
      7'o54: vJlF3gash = 32'd11698 ^ 32'b00000000000000000011111111111000 ^ 32'd4682;
      7'd100: vJlF3gash = 32'h7eba ^ 32'h7ebb;
      7'd94: vJlF3gash = 32'b00000000000000000010111011010111 ^ 32'b00000000000000000010111011010110;
      7'd37: vJlF3gash = 32'b00000000000000000011001111010010 ^ 32'b00000000000000000011001111010010;
      7'b0111101: vJlF3gash = 32'd8038 ^ 32'o17546;
      7'b1110010: vJlF3gash = 32'b00000000000000000100100001111101 ^ 32'h487c;
      7'b0111011: vJlF3gash = 32'd8561 ^ 32'd8560;
      7'd92: vJlF3gash = 32'b00000000000000000101101011011110 ^ 32'd23263;
      7'd4: vJlF3gash = 32'o22142 ^ 32'd25767 ^ 32'b00000000000000000100000011000101;
      7'd89: vJlF3gash = 32'b00000000000000000011001011101100 ^ 32'd15865 ^ 32'o7424;
      7'b1110110: vJlF3gash = 32'd6763 ^ 32'o15152;
      7'b1000000: vJlF3gash = 32'd7516 ^ 32'd19132 ^ 32'o53741;
      7'b1010110: vJlF3gash = 32'hafb ^ 32'hafa;
      7'hd: vJlF3gash = 32'o71073 ^ 32'h6441 ^ 32'h167a;
      7'h5f: vJlF3gash = 32'b00000000000000000101100011010011 ^ 32'o54322;
      7'b1111100: vJlF3gash = 32'h4052 ^ 32'b00000000000000000111011010011001 ^ 32'd14026;
      7'd35: vJlF3gash = 32'd24537 ^ 32'o40136 ^ 32'o17606;
      7'd122: vJlF3gash = 32'b00000000000000000110110001011001 ^ 32'o65410 ^ 32'o3520;
    endcase
  end

  logic [31:0] qaz6wx1C86;

  always_ff @(posedge clk_i) begin
    if(zZF) begin
      busy <= '0;
    end else begin
      busy <= vJlF3gash[32'b00000000000000000110010010101011 ^ 32'd21989 ^ 32'o30516];
    end
  end

  logic [31:0] q5Upj3TRGS8nkfV;
  always_comb begin
    case ({wKSnwVGWV, VICULOkZm, valid, eY8BfVPWv, XJhsywc8r, r0UH06pov5})
      6'd57: qaz6wx1C86 = 32'b00000000000000000100110110100011 ^ 32'd5756 ^ 32'b00000000000000000101101111011110;
      6'o32: qaz6wx1C86 = 32'h122b ^ 32'o35305 ^ 32'd10478;
      6'o70: qaz6wx1C86 = 32'h23a6 ^ 32'd9126;
      6'h17: qaz6wx1C86 = 32'b00000000000000000001010000110110 ^ 32'o64555 ^ 32'b00000000000000000111110101011011;
      6'd48: qaz6wx1C86 = 32'b00000000000000000111111111001010 ^ 32'b00000000000000000001011011100010 ^ 32'h6928;
      6'b100010: qaz6wx1C86 = 32'b00000000000000000011011000000111 ^ 32'd29847 ^ 32'b00000000000000000100001010010000;
      6'b101000: qaz6wx1C86 = 32'h5eb ^ 32'h5eb;
      6'o34: qaz6wx1C86 = 32'b00000000000000000001000000100001 ^ 32'o6036 ^ 32'd7231;
      6'd17: qaz6wx1C86 = 32'h4453 ^ 32'o35453 ^ 32'o77570;
      6'h3b: qaz6wx1C86 = 32'h4b98 ^ 32'b00000000000000000110011111010100 ^ 32'b00000000000000000010110001001100;
      6'o25: qaz6wx1C86 = 32'h1641 ^ 32'o14024 ^ 32'b00000000000000000000111001010101;
      6'o44: qaz6wx1C86 = 32'd13309 ^ 32'b00000000000000000100010111110000 ^ 32'b00000000000000000111011000001101;
      6'h27: qaz6wx1C86 = 32'o30762 ^ 32'b00000000000000000001011101001000 ^ 32'b00000000000000000010011010111011;
      6'o41: qaz6wx1C86 = 32'd3083 ^ 32'b00000000000000000000110000001010;
      6'o23: qaz6wx1C86 = 32'b00000000000000000100001001001000 ^ 32'hc84 ^ 32'o47314;
      6'd29: qaz6wx1C86 = 32'b00000000000000000011101000011101 ^ 32'b00000000000000000011101000011101;
      6'd32: qaz6wx1C86 = 32'd25103 ^ 32'o64407 ^ 32'hb08;
      6'o74: qaz6wx1C86 = 32'o72624 ^ 32'h7594;
      6'b101001: qaz6wx1C86 = 32'd12263 ^ 32'b00000000000000000110100010100001 ^ 32'b00000000000000000100011101000111;
      6'o17: qaz6wx1C86 = 32'd28762 ^ 32'o70132;
      6'd53: qaz6wx1C86 = 32'b00000000000000000111101110110101 ^ 32'b00000000000000000011100110010011 ^ 32'o41047;
      6'h10: qaz6wx1C86 = 32'd6743 ^ 32'o15127;
      6'b000100: qaz6wx1C86 = 32'd9356 ^ 32'd24233 ^ 32'o75045;
      6'b010100: qaz6wx1C86 = 32'h6c45 ^ 32'o66105;
      6'b111111: qaz6wx1C86 = 32'o16606 ^ 32'd17597 ^ 32'h593b;
      6'd42: qaz6wx1C86 = 32'o54744 ^ 32'd23012;
      6'b011000: qaz6wx1C86 = 32'o37063 ^ 32'b00000000000000000011111000110011;
      6'b101111: qaz6wx1C86 = 32'b00000000000000000101010111001110 ^ 32'd21967;
      6'b111110: qaz6wx1C86 = 32'b00000000000000000100100110001101 ^ 32'b00000000000000000011100100101101 ^ 32'd28832;
      6'o62: qaz6wx1C86 = 32'h7dc0 ^ 32'b00000000000000000110100000111010 ^ 32'h15fa;
      6'o53: qaz6wx1C86 = 32'b00000000000000000000001111100000 ^ 32'd29745 ^ 32'h77d0;
      6'o16: qaz6wx1C86 = 32'd7265 ^ 32'd7265;
      6'b011111: qaz6wx1C86 = 32'd14354 ^ 32'h3812;
      6'h9: qaz6wx1C86 = 32'b00000000000000000010000001110111 ^ 32'd8311;
      6'b100101: qaz6wx1C86 = 32'd24057 ^ 32'o5670 ^ 32'o53100;
      6'h1: qaz6wx1C86 = 32'h7c9b ^ 32'b00000000000000000111110010011011;
      6'h12: qaz6wx1C86 = 32'h6e4f ^ 32'd28239;
      6'o66: qaz6wx1C86 = 32'h4fae ^ 32'd17699 ^ 32'b00000000000000000000101010001101;
      6'o2: qaz6wx1C86 = 32'h5094 ^ 32'h5094;
      6'h8: qaz6wx1C86 = 32'd30330 ^ 32'h3b92 ^ 32'b00000000000000000100110111101000;
      6'd51: qaz6wx1C86 = 32'd10172 ^ 32'd10172;
      6'b101100: qaz6wx1C86 = 32'o26734 ^ 32'b00000000000000000011100111111001 ^ 32'd5157;
      6'h34: qaz6wx1C86 = 32'b00000000000000000101000110111000 ^ 32'd29643 ^ 32'b00000000000000000010001001110011;
      6'd55: qaz6wx1C86 = 32'h79aa ^ 32'h79aa;
      6'b010110: qaz6wx1C86 = 32'h403d ^ 32'h403d;
      6'b111101: qaz6wx1C86 = 32'd8081 ^ 32'h7365 ^ 32'h6cf5;
      6'd27: qaz6wx1C86 = 32'd26148 ^ 32'b00000000000000000100011001010110 ^ 32'h2072;
      6'h7: qaz6wx1C86 = 32'o46176 ^ 32'h4c7e;
      6'h2e: qaz6wx1C86 = 32'b00000000000000000010101111010010 ^ 32'd11218;
      6'o5: qaz6wx1C86 = 32'o47211 ^ 32'b00000000000000000100111010001001;
      6'o55: qaz6wx1C86 = 32'h1d5 ^ 32'd17801 ^ 32'h445d;
      6'b000110: qaz6wx1C86 = 32'b00000000000000000111100010000101 ^ 32'o65071 ^ 32'b00000000000000000001001010111100;
      6'd25: qaz6wx1C86 = 32'o64057 ^ 32'o64057;
      6'd11: qaz6wx1C86 = 32'b00000000000000000001111001101100 ^ 32'o17154;
      6'o72: qaz6wx1C86 = 32'o20634 ^ 32'h220c ^ 32'h390;
      6'd35: qaz6wx1C86 = 32'o60004 ^ 32'o35137 ^ 32'o55132;
      6'h3: qaz6wx1C86 = 32'h7a90 ^ 32'o14341 ^ 32'b00000000000000000110001001110001;
      6'h0: qaz6wx1C86 = 32'h529e ^ 32'b00000000000000000101001010011110;
      6'o14: qaz6wx1C86 = 32'h4869 ^ 32'o14172 ^ 32'h5013;
      6'd49: qaz6wx1C86 = 32'b00000000000000000101001111000011 ^ 32'h53c2;
      6'o12: qaz6wx1C86 = 32'b00000000000000000100101001110011 ^ 32'b00000000000000000100101001110011;
      6'b100110: qaz6wx1C86 = 32'h7f6 ^ 32'b00000000000000000000011111110110;
      6'd13: qaz6wx1C86 = 32'd29285 ^ 32'h5e43 ^ 32'd11302;
      6'b011110: qaz6wx1C86 = 32'o62031 ^ 32'b00000000000000000001011110101110 ^ 32'h73b7;
    endcase
  end

  assign r0UH06pov5 = UmLX == (32'o32572 ^ 32'h357a);

  always_ff @(posedge clk_i) begin
    if(zZF) begin
      valid <= '0;
    end else begin
      valid <= qaz6wx1C86[32'o46742 ^ 32'o24471 ^ 32'h64db];
    end
  end

  logic VVZKlkqbq;
  assign VVZKlkqbq = UmLX == (32'h73e2 ^ 32'b00000000000000000001101001001000 ^ 32'o64652);
  always_comb begin
    case ({wKSnwVGWV, VICULOkZm, VVZKlkqbq, XJhsywc8r})
      4'b1101: q5Upj3TRGS8nkfV = 32'h5ea0 ^ 32'hed25493;
      4'd3: q5Upj3TRGS8nkfV = 32'd15044 ^ 32'h3f17 ^ 32'b01011110010110011010111010001111;
      4'h6: q5Upj3TRGS8nkfV = 32'o34271 ^ 32'd4207 ^ 32'd832212430;
      4'o13: q5Upj3TRGS8nkfV = 32'o5247 ^ 32'h6d58 ^ 32'h6f961b2b;
      4'h0: q5Upj3TRGS8nkfV = 32'b00000000000000000001001011010010 ^ 32'o14336040213;
      4'd7: q5Upj3TRGS8nkfV = 32'd25270 ^ 32'h1bc519ae;
      4'o4: q5Upj3TRGS8nkfV = 32'd25792 ^ 32'b01010100100001001010111011011101;
      4'ha: q5Upj3TRGS8nkfV = 32'h60ab ^ 32'b00011110001100100000110100000110;
      4'hc: q5Upj3TRGS8nkfV = 32'h34a4 ^ 32'd13088 ^ 32'd102164953;
      4'o2: q5Upj3TRGS8nkfV = 32'b00000000000000000001000011001000 ^ 32'd1470131080;
      4'd5: q5Upj3TRGS8nkfV = 32'd3773 ^ 32'o14677436470;
      4'o17: q5Upj3TRGS8nkfV = 32'o31231 ^ 32'b01100100111110100100110000011011;
      4'b0001: q5Upj3TRGS8nkfV = 32'o36317 ^ 32'h6dbe ^ 32'b01010001100000101111011101101001;
      4'h8: q5Upj3TRGS8nkfV = 32'd3250 ^ 32'h1c00 ^ 32'h42d7eb62;
      4'b1110: q5Upj3TRGS8nkfV = 32'd2205 ^ 32'h3eb1 ^ 32'h74c58ad8;
      4'd9: q5Upj3TRGS8nkfV = 32'd13999 ^ 32'd25032 ^ 32'd1908358519;
    endcase
  end

  logic [31:0] eBnHjxu3POlmkT7;
  assign XJhsywc8r = FFDK4sD9m7 == (32'o26420 ^ 32'b00000000000000000011010010011010 ^ 32'h198b);
  always_comb begin
    case ({wKSnwVGWV, VICULOkZm, VVZKlkqbq, XJhsywc8r})
      4'd13: eBnHjxu3POlmkT7 = 32'o62772 ^ 32'd25234 ^ 32'd619253058;
      4'h9: eBnHjxu3POlmkT7 = 32'o37011 ^ 32'h78b64f90;
      4'h5: eBnHjxu3POlmkT7 = 32'd5655 ^ 32'd13393 ^ 32'o14774560176;
      4'b0011: eBnHjxu3POlmkT7 = 32'h421e ^ 32'o24300 ^ 32'h33beeb7f;
      4'b1110: eBnHjxu3POlmkT7 = 32'hff7 ^ 32'b00000000000000000010100001011010 ^ 32'b01111101110010100011111011111010;
      4'h7: eBnHjxu3POlmkT7 = 32'o65020 ^ 32'o16034426322;
      4'b0100: eBnHjxu3POlmkT7 = 32'h6c1b ^ 32'd1616384739;
      4'd15: eBnHjxu3POlmkT7 = 32'b00000000000000000011100111110011 ^ 32'h6d8d37c6;
      4'h2: eBnHjxu3POlmkT7 = 32'o14042 ^ 32'd25336 ^ 32'o2654636133;
      4'b0110: eBnHjxu3POlmkT7 = 32'b00000000000000000100000000010100 ^ 32'o75031 ^ 32'h1a1b1874;
      4'b0001: eBnHjxu3POlmkT7 = 32'b00000000000000000100010000101001 ^ 32'b00000000000000000101011101101000 ^ 32'h2ef4b8b3;
      4'd8: eBnHjxu3POlmkT7 = 32'h140c ^ 32'b00000000000000000000010110101001 ^ 32'b01101100000110101011001000011111;
      4'hb: eBnHjxu3POlmkT7 = 32'b00000000000000000001001000000010 ^ 32'b00000000000000000101011100000010 ^ 32'b00101111110001001001110111011101;
      4'b1010: eBnHjxu3POlmkT7 = 32'o64005 ^ 32'd1843325073;
      4'h0: eBnHjxu3POlmkT7 = 32'h1a2d ^ 32'd734609828;
      4'd12: eBnHjxu3POlmkT7 = 32'b00000000000000000011101111111110 ^ 32'b01110001100110001001111110011100;
    endcase
  end

  always_ff @(posedge clk_i) begin
    if(zZF) begin
      data <= '0;
    end else if (q5Upj3TRGS8nkfV[32'd23241 ^ 32'b00000000000000000101101011001000]) begin
      data <= '0;
    end else if(eBnHjxu3POlmkT7[32'o72553 ^ 32'b00000000000000000111010101101001]) begin
      data <= FFDK4sD9m7;
    end
    else begin
      data <= data;
    end
  end

  assign fcS5S0IailtPh = UmLX == (32'o13330 ^ 32'o43045 ^ 32'd20721);
  logic [31:0] SuhrzWcGiwP2SmTaYCK;
  always_comb begin
    case ({wKSnwVGWV, fcS5S0IailtPh, VICULOkZm, XJhsywc8r})
      4'd5: SuhrzWcGiwP2SmTaYCK = 32'h664e ^ 32'o31120 ^ 32'h121a79bb;
      4'h4: SuhrzWcGiwP2SmTaYCK = 32'h3c52 ^ 32'o16325204045;
      4'h1: SuhrzWcGiwP2SmTaYCK = 32'd15965 ^ 32'd2111526847;
      4'd13: SuhrzWcGiwP2SmTaYCK = 32'd13874 ^ 32'b00000000000000000110000010010010 ^ 32'b01111110111010011111001101110001;
      4'd8: SuhrzWcGiwP2SmTaYCK = 32'b00000000000000000110010001000100 ^ 32'o1651 ^ 32'h39cc7d3b;
      4'hc: SuhrzWcGiwP2SmTaYCK = 32'o6065 ^ 32'd343741462;
      4'b1011: SuhrzWcGiwP2SmTaYCK = 32'h6239 ^ 32'h5501 ^ 32'o6775127066;
      4'd10: SuhrzWcGiwP2SmTaYCK = 32'o34075 ^ 32'o6174646137;
      4'd3: SuhrzWcGiwP2SmTaYCK = 32'b00000000000000000001001001010110 ^ 32'h26c0 ^ 32'd368251297;
      4'd2: SuhrzWcGiwP2SmTaYCK = 32'h6859 ^ 32'b00000110101101000010000000111010;
      4'o7: SuhrzWcGiwP2SmTaYCK = 32'h3a47 ^ 32'd1161903040;
      4'he: SuhrzWcGiwP2SmTaYCK = 32'b00000000000000000000101000101011 ^ 32'o17563345053;
      4'h9: SuhrzWcGiwP2SmTaYCK = 32'o7100 ^ 32'o15764422501;
      4'o6: SuhrzWcGiwP2SmTaYCK = 32'd4171 ^ 32'd30744 ^ 32'd6904852;
      4'd15: SuhrzWcGiwP2SmTaYCK = 32'o32047 ^ 32'o30752 ^ 32'b01110010010101100100010111100000;
      4'd0: SuhrzWcGiwP2SmTaYCK = 32'h1460 ^ 32'h5567 ^ 32'd882296647;
    endcase
  end

  logic [31:0] FHGBch0qBHxqcbX8Dlb;
  always_comb begin
    case ({wKSnwVGWV, fcS5S0IailtPh, VICULOkZm, XJhsywc8r})
      4'd12: FHGBch0qBHxqcbX8Dlb = 32'b00000000000000000000110001001011 ^ 32'h331f09ba;
      4'd15: FHGBch0qBHxqcbX8Dlb = 32'd2624 ^ 32'b00111010001111100110100101010111;
      4'd0: FHGBch0qBHxqcbX8Dlb = 32'h6a79 ^ 32'o11016714577;
      4'h4: FHGBch0qBHxqcbX8Dlb = 32'o36147 ^ 32'b00000110001011010101001100101101;
      4'd14: FHGBch0qBHxqcbX8Dlb = 32'd24643 ^ 32'h635a ^ 32'h36813882;
      4'ha: FHGBch0qBHxqcbX8Dlb = 32'b00000000000000000011100001010010 ^ 32'b00000000000000000100110000111010 ^ 32'o2211317713;
      4'b1011: FHGBch0qBHxqcbX8Dlb = 32'o61116 ^ 32'h1202 ^ 32'h21745a02;
      4'o2: FHGBch0qBHxqcbX8Dlb = 32'd26734 ^ 32'o16770 ^ 32'h4fc6d1d5;
      4'b0101: FHGBch0qBHxqcbX8Dlb = 32'o63144 ^ 32'o67521 ^ 32'h714246f3;
      4'b0110: FHGBch0qBHxqcbX8Dlb = 32'o10140 ^ 32'h427bb924;
      4'h1: FHGBch0qBHxqcbX8Dlb = 32'o12166 ^ 32'h1268 ^ 32'b01101001010000011001010010110110;
      4'd13: FHGBch0qBHxqcbX8Dlb = 32'h3647 ^ 32'o16622 ^ 32'b01110110001010000111000100101100;
      4'h9: FHGBch0qBHxqcbX8Dlb = 32'b00000000000000000000111001010101 ^ 32'b01001011011110100011011100111100;
      4'h7: FHGBch0qBHxqcbX8Dlb = 32'o35134 ^ 32'h459eecf4;
      4'h8: FHGBch0qBHxqcbX8Dlb = 32'd25689 ^ 32'o40251 ^ 32'h3a6f4fd0;
      4'o3: FHGBch0qBHxqcbX8Dlb = 32'd4715 ^ 32'h63c1 ^ 32'b01001111110001011111010111000100;
    endcase
  end

  always_ff @(posedge clk_i) begin
    if(zZF) begin
      baudrate <= '0;
    end else if (SuhrzWcGiwP2SmTaYCK[32'd3188 ^ 32'b00000000000000000000110001110111]) begin
      baudrate <= '0;
    end
    else if(FHGBch0qBHxqcbX8Dlb[32'b00000000000000000000110101101111 ^ 32'h787d ^ 32'o72426]) begin
      baudrate <= FFDK4sD9m7;
    end
    else begin
      baudrate <= baudrate;
    end
  end

  logic [31:0] WLGbSSV5YzHmlpmqLI;

  logic [31:0] b5l5UfftZRDTX1AD2;
  logic m4Js9aFV4Us;
  always_comb begin
    case ({wKSnwVGWV, m4Js9aFV4Us, VICULOkZm, XJhsywc8r})
      4'd14: b5l5UfftZRDTX1AD2 = 32'b00000000000000000110010110000000 ^ 32'd295811877;
      4'b0111: b5l5UfftZRDTX1AD2 = 32'h159d ^ 32'o12602005631;
      4'd6: b5l5UfftZRDTX1AD2 = 32'h6ba0 ^ 32'o11557450265;
      4'd2: b5l5UfftZRDTX1AD2 = 32'h43af ^ 32'd17152 ^ 32'h22f4f996;
      4'b1101: b5l5UfftZRDTX1AD2 = 32'b00000000000000000011101110000100 ^ 32'h1e89d3c;
      4'o13: b5l5UfftZRDTX1AD2 = 32'o63613 ^ 32'o15557237564;
      4'd1: b5l5UfftZRDTX1AD2 = 32'd6578 ^ 32'o2423507117;
      4'b1111: b5l5UfftZRDTX1AD2 = 32'b00000000000000000000111101111101 ^ 32'd5106 ^ 32'b00101010110111011010011011110000;
      4'h4: b5l5UfftZRDTX1AD2 = 32'h17a8 ^ 32'd1199459581;
      4'o5: b5l5UfftZRDTX1AD2 = 32'b00000000000000000100000110100100 ^ 32'b00000000000000000001010001011000 ^ 32'h2acd6c79;
      4'd3: b5l5UfftZRDTX1AD2 = 32'h6dab ^ 32'd2104322542;
      4'o10: b5l5UfftZRDTX1AD2 = 32'o64626 ^ 32'd407919674;
      4'b1100: b5l5UfftZRDTX1AD2 = 32'h1187 ^ 32'd17050 ^ 32'b00100101100100001010000100001000;
      4'h9: b5l5UfftZRDTX1AD2 = 32'd5010 ^ 32'd28993 ^ 32'b01000000000011010011100101100111;
      4'b0000: b5l5UfftZRDTX1AD2 = 32'o67666 ^ 32'o33557 ^ 32'd1228297272;
      4'o12: b5l5UfftZRDTX1AD2 = 32'b00000000000000000011110110001110 ^ 32'b00000000000000000011011100001001 ^ 32'o15300071342;
    endcase
  end

  logic [31:0] fhHTYz8JNP73GgkZp;
  always_comb begin
    case ({wKSnwVGWV, m4Js9aFV4Us, VICULOkZm, XJhsywc8r})
      4'd6: fhHTYz8JNP73GgkZp = 32'o47241 ^ 32'o62175 ^ 32'd458013848;
      4'ha: fhHTYz8JNP73GgkZp = 32'b00000000000000000111011010010011 ^ 32'b00110011011111001110001010000110;
      4'o7: fhHTYz8JNP73GgkZp = 32'b00000000000000000111100010011110 ^ 32'h7dcc2c86;
      4'o10: fhHTYz8JNP73GgkZp = 32'h229a ^ 32'b00000000000000000111000000001110 ^ 32'h1202b248;
      4'o13: fhHTYz8JNP73GgkZp = 32'b00000000000000000010000010001111 ^ 32'b00000000000000000100000101100110 ^ 32'o13251517010;
      4'b0000: fhHTYz8JNP73GgkZp = 32'o51267 ^ 32'b00000000000000000100000111001100 ^ 32'd110940771;
      4'd1: fhHTYz8JNP73GgkZp = 32'o76263 ^ 32'h3675cebe;
      4'h4: fhHTYz8JNP73GgkZp = 32'o75250 ^ 32'b00011100000101100010111010111001;
      4'b1110: fhHTYz8JNP73GgkZp = 32'd18561 ^ 32'd1483794795;
      4'h9: fhHTYz8JNP73GgkZp = 32'd19606 ^ 32'o32726 ^ 32'd980015896;
      4'o3: fhHTYz8JNP73GgkZp = 32'd20652 ^ 32'b00000000000000000001001100100101 ^ 32'd868638757;
      4'h2: fhHTYz8JNP73GgkZp = 32'o23260 ^ 32'h19035575;
      4'hd: fhHTYz8JNP73GgkZp = 32'd7812 ^ 32'b00000000000000000001001010111111 ^ 32'o16052401775;
      4'b1100: fhHTYz8JNP73GgkZp = 32'b00000000000000000100101010001100 ^ 32'o13236356763;
      4'o5: fhHTYz8JNP73GgkZp = 32'o22245 ^ 32'b00000111001111101010111000101001;
      4'o17: fhHTYz8JNP73GgkZp = 32'b00000000000000000111001001111101 ^ 32'd7759 ^ 32'b00100111001011110111011100110001;
    endcase
  end
  assign m4Js9aFV4Us = UmLX == (32'd22117 ^ 32'd32555 ^ 32'd10590);

  always_ff @(posedge clk_i) begin
    if(zZF) begin
      parity_en <= '0;
    end else if (b5l5UfftZRDTX1AD2[32'h7906 ^ 32'h12c0 ^ 32'h6bc7]) begin
      parity_en <= '0;
    end
    else if(fhHTYz8JNP73GgkZp[32'o1770 ^ 32'o1771]) begin
      parity_en <= FFDK4sD9m7;
    end
    else begin
      parity_en <= parity_en;
    end
  end

  logic P0EEllcI4VCU;
  assign P0EEllcI4VCU = UmLX == (32'o62726 ^ 32'd26050);
  always_comb begin
    case ({m4Js9aFV4Us, P0EEllcI4VCU, VICULOkZm, XJhsywc8r, wKSnwVGWV, fcS5S0IailtPh})
      6'b010011: WLGbSSV5YzHmlpmqLI = 32'h7a7f ^ 32'o6421703407;
      6'h1a: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000100101001100010 ^ 32'h62321c5f;
      6'h2f: WLGbSSV5YzHmlpmqLI = 32'o63023 ^ 32'h722d90fd;
      6'd28: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000001111001011011 ^ 32'h3d02 ^ 32'd1738296917;
      6'he: WLGbSSV5YzHmlpmqLI = 32'd10385 ^ 32'h1e9099e6;
      6'b000110: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000010111010110001 ^ 32'd100341241;
      6'h7: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000101100010101101 ^ 32'o74006 ^ 32'h4af4ca7f;
      6'd53: WLGbSSV5YzHmlpmqLI = 32'h61fd ^ 32'd21334 ^ 32'b01101010110001001001010101000010;
      6'o61: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000011101000001100 ^ 32'd1070093101;
      6'o76: WLGbSSV5YzHmlpmqLI = 32'h5d9 ^ 32'o4453034147;
      6'd36: WLGbSSV5YzHmlpmqLI = 32'o67076 ^ 32'o65503 ^ 32'o236115274;
      6'h29: WLGbSSV5YzHmlpmqLI = 32'o40054 ^ 32'b00000000000000000100100000101100 ^ 32'd438005057;
      6'b111011: WLGbSSV5YzHmlpmqLI = 32'h7e4 ^ 32'h5a9eb098;
      6'o21: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000010011010000110 ^ 32'o73640 ^ 32'b00101111111101010100111111100010;
      6'd40: WLGbSSV5YzHmlpmqLI = 32'h1630 ^ 32'b01100011100010011101000101001101;
      6'h37: WLGbSSV5YzHmlpmqLI = 32'd13814 ^ 32'd1499541943;
      6'o17: WLGbSSV5YzHmlpmqLI = 32'h528d ^ 32'h6c10 ^ 32'o7462474716;
      6'd34: WLGbSSV5YzHmlpmqLI = 32'd6725 ^ 32'b01111010100000111001101011110101;
      6'd2: WLGbSSV5YzHmlpmqLI = 32'o3277 ^ 32'h1b1d ^ 32'd1165033499;
      6'h30: WLGbSSV5YzHmlpmqLI = 32'h100f ^ 32'b00000000000000000111011001101110 ^ 32'o6552062231;
      6'b010110: WLGbSSV5YzHmlpmqLI = 32'o74164 ^ 32'd1434393388;
      6'b111101: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000101101111011101 ^ 32'b00000000000000000100011101100000 ^ 32'd909162724;
      6'd57: WLGbSSV5YzHmlpmqLI = 32'd2543 ^ 32'b00001000011000100101001011101011;
      6'b101011: WLGbSSV5YzHmlpmqLI = 32'd15905 ^ 32'o14605 ^ 32'd426889412;
      6'o72: WLGbSSV5YzHmlpmqLI = 32'd13291 ^ 32'o13620560216;
      6'b011111: WLGbSSV5YzHmlpmqLI = 32'd7248 ^ 32'h39d2009f;
      6'b101100: WLGbSSV5YzHmlpmqLI = 32'o64036 ^ 32'd2115225742;
      6'o46: WLGbSSV5YzHmlpmqLI = 32'd16951 ^ 32'b00000000000000000111011011010100 ^ 32'b01011100001111100101001100110011;
      6'b100011: WLGbSSV5YzHmlpmqLI = 32'o42102 ^ 32'b00000000000000000010010101111011 ^ 32'b01100001010001000101101011010101;
      6'o30: WLGbSSV5YzHmlpmqLI = 32'o46155 ^ 32'b00001111100010110010101101111001;
      6'h12: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000101000010000010 ^ 32'h3d68 ^ 32'o5006130516;
      6'o52: WLGbSSV5YzHmlpmqLI = 32'h1425 ^ 32'd21437 ^ 32'h6c10c5c1;
      6'o35: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000100100001010111 ^ 32'b00001111100001110110000101101011;
      6'd13: WLGbSSV5YzHmlpmqLI = 32'd32404 ^ 32'o5267624761;
      6'b111000: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000101111111110011 ^ 32'd9391 ^ 32'b00000010001110111100111110000100;
      6'd63: WLGbSSV5YzHmlpmqLI = 32'o27726 ^ 32'd21232 ^ 32'h60c73c71;
      6'b100111: WLGbSSV5YzHmlpmqLI = 32'h6c33 ^ 32'd1348383130;
      6'h33: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000000111000000101 ^ 32'b00000000000000000100011111000110 ^ 32'o1413653112;
      6'b110010: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000110010000001000 ^ 32'b00101000100110011110100011100100;
      6'h8: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000010110010100110 ^ 32'o11036124126;
      6'b100000: WLGbSSV5YzHmlpmqLI = 32'd17996 ^ 32'd55914332;
      6'o3: WLGbSSV5YzHmlpmqLI = 32'o30274 ^ 32'o4415063561;
      6'o11: WLGbSSV5YzHmlpmqLI = 32'h56a3 ^ 32'o44537 ^ 32'o7406347521;
      6'o13: WLGbSSV5YzHmlpmqLI = 32'd10907 ^ 32'd1539340531;
      6'h25: WLGbSSV5YzHmlpmqLI = 32'h183a ^ 32'h321abce3;
      6'b110110: WLGbSSV5YzHmlpmqLI = 32'hbfa ^ 32'b00000000000000000001100100011111 ^ 32'o13474325645;
      6'h17: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000010001001110000 ^ 32'o15121 ^ 32'd1851010648;
      6'b001100: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000101010010011000 ^ 32'h1ab7 ^ 32'o2022343312;
      6'o36: WLGbSSV5YzHmlpmqLI = 32'o71124 ^ 32'o44222 ^ 32'o7444464371;
      6'd46: WLGbSSV5YzHmlpmqLI = 32'o36027 ^ 32'o65335 ^ 32'd371448084;
      6'b010000: WLGbSSV5YzHmlpmqLI = 32'h7c89 ^ 32'd1941236341;
      6'b010100: WLGbSSV5YzHmlpmqLI = 32'h247b ^ 32'o44370 ^ 32'd1196722951;
      6'd27: WLGbSSV5YzHmlpmqLI = 32'd29790 ^ 32'o73472 ^ 32'h5602858c;
      6'b000101: WLGbSSV5YzHmlpmqLI = 32'd1205 ^ 32'h6c76 ^ 32'd1912730239;
      6'b011001: WLGbSSV5YzHmlpmqLI = 32'h2066 ^ 32'h6ba9 ^ 32'd942376155;
      6'o1: WLGbSSV5YzHmlpmqLI = 32'o56303 ^ 32'b00111110001100010100011111001011;
      6'o4: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000101101010111000 ^ 32'h4fc2c804;
      6'h34: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000011100000000001 ^ 32'o13201041555;
      6'd45: WLGbSSV5YzHmlpmqLI = 32'b00000000000000000001001000011010 ^ 32'b00000000000000000010010100010101 ^ 32'hb1fbcbe;
      6'b001010: WLGbSSV5YzHmlpmqLI = 32'd159 ^ 32'd1516813251;
      6'b010101: WLGbSSV5YzHmlpmqLI = 32'o47170 ^ 32'h693d2bc0;
      6'd60: WLGbSSV5YzHmlpmqLI = 32'h31e1 ^ 32'd1326516696;
      6'h21: WLGbSSV5YzHmlpmqLI = 32'd28745 ^ 32'o14753 ^ 32'o102622513;
      6'h0: WLGbSSV5YzHmlpmqLI = 32'd12999 ^ 32'd3981 ^ 32'o16012611657;
    endcase
  end

  assign wKSnwVGWV  = pEo &  qICjuvAOmWmr;
  assign VICULOkZm = UmLX == (32'h148f ^ 32'o12253);

  logic [31:0] vBjc8EzRDlz48WXa4k;
  always_comb begin
    case ({m4Js9aFV4Us, P0EEllcI4VCU, VICULOkZm, XJhsywc8r, wKSnwVGWV, fcS5S0IailtPh})
      6'd9: vBjc8EzRDlz48WXa4k = 32'b00000000000000000001110000100110 ^ 32'd1968865001;
      6'b110111: vBjc8EzRDlz48WXa4k = 32'b00000000000000000111101101111010 ^ 32'b00000000000000000100111000100110 ^ 32'o10303624447;
      6'h38: vBjc8EzRDlz48WXa4k = 32'o47563 ^ 32'd22966 ^ 32'b01011000111000010111000111010011;
      6'b001110: vBjc8EzRDlz48WXa4k = 32'd28180 ^ 32'd1770718541;
      6'd44: vBjc8EzRDlz48WXa4k = 32'o26641 ^ 32'o47214 ^ 32'd1269075633;
      6'b101101: vBjc8EzRDlz48WXa4k = 32'h579e ^ 32'o6642351503;
      6'o76: vBjc8EzRDlz48WXa4k = 32'h4b5d ^ 32'b00000000000000000111110001100111 ^ 32'd2002868800;
      6'o31: vBjc8EzRDlz48WXa4k = 32'd26089 ^ 32'b00000000000000000101101011101001 ^ 32'h25c93bcb;
      6'd30: vBjc8EzRDlz48WXa4k = 32'b00000000000000000011011111010111 ^ 32'h4bcd7ab8;
      6'h3f: vBjc8EzRDlz48WXa4k = 32'h755a ^ 32'h683eb3f6;
      6'd50: vBjc8EzRDlz48WXa4k = 32'o24614 ^ 32'o741700252;
      6'b110001: vBjc8EzRDlz48WXa4k = 32'b00000000000000000111111110001111 ^ 32'b00000000000000000010101101110101 ^ 32'h25a4e761;
      6'b101011: vBjc8EzRDlz48WXa4k = 32'b00000000000000000000001110100101 ^ 32'd2244 ^ 32'h68c578ae;
      6'h5: vBjc8EzRDlz48WXa4k = 32'b00000000000000000111010000110101 ^ 32'h217d ^ 32'd278675848;
      6'o60: vBjc8EzRDlz48WXa4k = 32'o52623 ^ 32'd1522064583;
      6'o17: vBjc8EzRDlz48WXa4k = 32'd6161 ^ 32'o55517 ^ 32'b01001001001111001110001011011010;
      6'o50: vBjc8EzRDlz48WXa4k = 32'd1456 ^ 32'h4076583a;
      6'o24: vBjc8EzRDlz48WXa4k = 32'h69ff ^ 32'd1647636143;
      6'o47: vBjc8EzRDlz48WXa4k = 32'd23475 ^ 32'o13355467573;
      6'o52: vBjc8EzRDlz48WXa4k = 32'h59a9 ^ 32'd269481827;
      6'o71: vBjc8EzRDlz48WXa4k = 32'd31087 ^ 32'h7630562;
      6'h18: vBjc8EzRDlz48WXa4k = 32'o35755 ^ 32'h6a83bd37;
      6'd29: vBjc8EzRDlz48WXa4k = 32'o6733 ^ 32'h4a379444;
      6'd7: vBjc8EzRDlz48WXa4k = 32'h482e ^ 32'o26415 ^ 32'h159216ab;
      6'd28: vBjc8EzRDlz48WXa4k = 32'o61737 ^ 32'o26101 ^ 32'h12fd684a;
      6'o22: vBjc8EzRDlz48WXa4k = 32'o13006 ^ 32'o26247 ^ 32'b01011001100101010111010000011010;
      6'o32: vBjc8EzRDlz48WXa4k = 32'd4070 ^ 32'h20b1 ^ 32'd1493582438;
      6'd8: vBjc8EzRDlz48WXa4k = 32'h722a ^ 32'd29398 ^ 32'd1335986429;
      6'd16: vBjc8EzRDlz48WXa4k = 32'b00000000000000000100001000001101 ^ 32'h2117 ^ 32'o7123071615;
      6'd0: vBjc8EzRDlz48WXa4k = 32'b00000000000000000111100001001010 ^ 32'h7ecc ^ 32'b00111101001001011100000000011001;
      6'd13: vBjc8EzRDlz48WXa4k = 32'h4418 ^ 32'h4fbe ^ 32'o10512704470;
      6'd46: vBjc8EzRDlz48WXa4k = 32'h19a ^ 32'b00000000000000000101101000011100 ^ 32'h50de6cc1;
      6'b100110: vBjc8EzRDlz48WXa4k = 32'd1979 ^ 32'b00101111001000100000011100100000;
      6'b101001: vBjc8EzRDlz48WXa4k = 32'h2fac ^ 32'o76464 ^ 32'd1859925953;
      6'h3: vBjc8EzRDlz48WXa4k = 32'o20074 ^ 32'd1241899107;
      6'o33: vBjc8EzRDlz48WXa4k = 32'o34742 ^ 32'b00001000000101001000010101000110;
      6'hc: vBjc8EzRDlz48WXa4k = 32'b00000000000000000001101000011100 ^ 32'o14507726611;
      6'd2: vBjc8EzRDlz48WXa4k = 32'h4c43 ^ 32'h5dfc9c0f;
      6'd51: vBjc8EzRDlz48WXa4k = 32'o51610 ^ 32'o2712712356;
      6'd61: vBjc8EzRDlz48WXa4k = 32'd8545 ^ 32'o5010064657;
      6'd52: vBjc8EzRDlz48WXa4k = 32'h7d85 ^ 32'b00000000000000000111110011001110 ^ 32'o2373371533;
      6'o23: vBjc8EzRDlz48WXa4k = 32'h4002 ^ 32'h7270 ^ 32'o13661424031;
      6'd47: vBjc8EzRDlz48WXa4k = 32'd11159 ^ 32'o17745 ^ 32'd1507346480;
      6'b001011: vBjc8EzRDlz48WXa4k = 32'b00000000000000000111000000011111 ^ 32'o16126427520;
      6'd34: vBjc8EzRDlz48WXa4k = 32'o57711 ^ 32'o47362 ^ 32'o6556706570;
      6'b010001: vBjc8EzRDlz48WXa4k = 32'd27658 ^ 32'o13440363525;
      6'd53: vBjc8EzRDlz48WXa4k = 32'b00000000000000000010011110000001 ^ 32'd923797700;
      6'h20: vBjc8EzRDlz48WXa4k = 32'b00000000000000000000101111010000 ^ 32'b00001111101110010101110100011011;
      6'o6: vBjc8EzRDlz48WXa4k = 32'o17061 ^ 32'o10271662043;
      6'o4: vBjc8EzRDlz48WXa4k = 32'o45070 ^ 32'b00010101110001010001001000101000;
      6'ha: vBjc8EzRDlz48WXa4k = 32'b00000000000000000100011000100011 ^ 32'o77146 ^ 32'o5725726402;
      6'h17: vBjc8EzRDlz48WXa4k = 32'o10761 ^ 32'o47530 ^ 32'd846604252;
      6'o37: vBjc8EzRDlz48WXa4k = 32'd25044 ^ 32'o76632 ^ 32'o12032654357;
      6'b111010: vBjc8EzRDlz48WXa4k = 32'd9068 ^ 32'd1215680840;
      6'o45: vBjc8EzRDlz48WXa4k = 32'd23998 ^ 32'o20113 ^ 32'o11606433661;
      6'o1: vBjc8EzRDlz48WXa4k = 32'o21107 ^ 32'd17556 ^ 32'o2065074715;
      6'b100100: vBjc8EzRDlz48WXa4k = 32'h33c2 ^ 32'b00000000000000000101101010000011 ^ 32'b00000110011010101111000010000000;
      6'o26: vBjc8EzRDlz48WXa4k = 32'h67f4 ^ 32'o14126711433;
      6'o25: vBjc8EzRDlz48WXa4k = 32'h3df8 ^ 32'b01011010011010110100011011110000;
      6'o43: vBjc8EzRDlz48WXa4k = 32'b00000000000000000000100111000101 ^ 32'h74b56408;
      6'o73: vBjc8EzRDlz48WXa4k = 32'b00000000000000000100110101101000 ^ 32'b00000000000000000010101100001111 ^ 32'b01110110100101111011001000011000;
      6'o66: vBjc8EzRDlz48WXa4k = 32'd20862 ^ 32'd2142 ^ 32'b01011110101000000011101011001001;
      6'd60: vBjc8EzRDlz48WXa4k = 32'd30564 ^ 32'b01100101011101001001000011101011;
      6'b100001: vBjc8EzRDlz48WXa4k = 32'b00000000000000000011010111001101 ^ 32'b00100101111010001111100000001000;
    endcase
  end

  logic [31:0] jMTaMbqs055c0zWDyuyX;
  always_comb begin
    case ({VICULOkZm, XJhsywc8r, wKSnwVGWV, pEo, qICjuvAOmWmr})
      5'ha: jMTaMbqs055c0zWDyuyX = 32'o73053 ^ 32'd2060447563;
      5'd1: jMTaMbqs055c0zWDyuyX = 32'd21071 ^ 32'b00001110111001010101111011000110;
      5'o36: jMTaMbqs055c0zWDyuyX = 32'o63740 ^ 32'h70d4 ^ 32'b01010001001001000110011110010010;
      5'o3: jMTaMbqs055c0zWDyuyX = 32'd9800 ^ 32'o4546566315;
      5'd23: jMTaMbqs055c0zWDyuyX = 32'b00000000000000000001011111111100 ^ 32'h4293 ^ 32'h38506077;
      5'h18: jMTaMbqs055c0zWDyuyX = 32'd16889 ^ 32'b01111111000001000101110000010000;
      5'h1f: jMTaMbqs055c0zWDyuyX = 32'h11dc ^ 32'h6066bf0e;
      5'hc: jMTaMbqs055c0zWDyuyX = 32'b00000000000000000100101000100100 ^ 32'd17145 ^ 32'b01111001101001110100010101100100;
      5'b10110: jMTaMbqs055c0zWDyuyX = 32'd28160 ^ 32'd1424638173;
      5'd17: jMTaMbqs055c0zWDyuyX = 32'd7186 ^ 32'h1fe2 ^ 32'h3f956080;
      5'b11010: jMTaMbqs055c0zWDyuyX = 32'h15f2 ^ 32'd5099 ^ 32'h4913b6d4;
      5'h9: jMTaMbqs055c0zWDyuyX = 32'h4c2f ^ 32'h71a0 ^ 32'b00001100000001010001000000000011;
      5'd29: jMTaMbqs055c0zWDyuyX = 32'h3de3 ^ 32'b00101001010010010101111101110110;
      5'o16: jMTaMbqs055c0zWDyuyX = 32'o17035 ^ 32'h4e89 ^ 32'h7bdf00ac;
      5'd15: jMTaMbqs055c0zWDyuyX = 32'h4819 ^ 32'd5201 ^ 32'b00110000101110111110101010011101;
      5'o4: jMTaMbqs055c0zWDyuyX = 32'd20548 ^ 32'h10344c94;
      5'b11001: jMTaMbqs055c0zWDyuyX = 32'o65765 ^ 32'o47043 ^ 32'b01100100111111110111000011100011;
      5'b00101: jMTaMbqs055c0zWDyuyX = 32'd31297 ^ 32'd5304 ^ 32'h23b36249;
      5'd19: jMTaMbqs055c0zWDyuyX = 32'b00000000000000000111000000001011 ^ 32'o4472612632;
      5'd2: jMTaMbqs055c0zWDyuyX = 32'b00000000000000000111110001001100 ^ 32'd17247 ^ 32'h555c1aef;
      5'd28: jMTaMbqs055c0zWDyuyX = 32'h13e7 ^ 32'b00010111110000011101010111100011;
      5'b10100: jMTaMbqs055c0zWDyuyX = 32'h1a07 ^ 32'h713a ^ 32'h7b647c68;
      5'd27: jMTaMbqs055c0zWDyuyX = 32'd27114 ^ 32'h1f7c ^ 32'b00111111111000011101110000111011;
      5'h6: jMTaMbqs055c0zWDyuyX = 32'h243d ^ 32'd484145837;
      5'd13: jMTaMbqs055c0zWDyuyX = 32'o72040 ^ 32'o6326065451;
      5'h7: jMTaMbqs055c0zWDyuyX = 32'b00000000000000000100111000111010 ^ 32'h2048 ^ 32'b00010100100110011101000001011011;
      5'h15: jMTaMbqs055c0zWDyuyX = 32'b00000000000000000100010000000100 ^ 32'h37ed0d9d;
      5'b10010: jMTaMbqs055c0zWDyuyX = 32'b00000000000000000100011000001110 ^ 32'd26026 ^ 32'd2088858357;
      5'o0: jMTaMbqs055c0zWDyuyX = 32'd10323 ^ 32'd460283331;
      5'hb: jMTaMbqs055c0zWDyuyX = 32'o20050 ^ 32'd438053772;
      5'o10: jMTaMbqs055c0zWDyuyX = 32'o74066 ^ 32'b00000000000000000110011000010000 ^ 32'o1737740073;
      5'b10000: jMTaMbqs055c0zWDyuyX = 32'b00000000000000000111001000010110 ^ 32'd212527463;
    endcase
  end

  logic [31:0] cI7ozekBmfu12;
  always_comb begin
    case ({VICULOkZm, XJhsywc8r, wKSnwVGWV, pEo, qICjuvAOmWmr})
      5'b01000: cI7ozekBmfu12 = 32'd290915043 ^ 32'o20660661050 ^ 32'hd1d90202;
      5'o31: cI7ozekBmfu12 = 32'd297552609 ^ 32'o11767541767;
      5'b00010: cI7ozekBmfu12 = 32'o5423064466 ^ 32'b00111011000010000111100010001101;
      5'h9: cI7ozekBmfu12 = 32'o4100311461 ^ 32'o7220423007 ^ 32'd903897080;
      5'h17: cI7ozekBmfu12 = 32'o23642451113 ^ 32'ha14628c7 ^ 32'b00101101000001110100000001010010;
      5'b00101: cI7ozekBmfu12 = 32'd3528236378 ^ 32'b10100011000110010010110001001011;
      5'h1f: cI7ozekBmfu12 = 32'hf6ab601a ^ 32'hd200c845;
      5'hd: cI7ozekBmfu12 = 32'o16770665634 ^ 32'd165392386 ^ 32'h6310ab4e;
      5'd6: cI7ozekBmfu12 = 32'hebb4c65 ^ 32'b00100000110011011111110000101110;
      5'o36: cI7ozekBmfu12 = 32'b10101111001011000000001011100010 ^ 32'o37573560442;
      5'h7: cI7ozekBmfu12 = 32'b10101001000000100011110000001010 ^ 32'hd51c6a98;
      5'b11000: cI7ozekBmfu12 = 32'd1232251627 ^ 32'o502717172 ^ 32'o203247034;
      5'b01100: cI7ozekBmfu12 = 32'o15575165117 ^ 32'b01100010011000111011001010000100;
      5'd21: cI7ozekBmfu12 = 32'd3119711741 ^ 32'd3765016980 ^ 32'o11466474470;
      5'b11101: cI7ozekBmfu12 = 32'b11011001100000111100100010101100 ^ 32'h4eafab5d ^ 32'd3050190571;
      5'b11011: cI7ozekBmfu12 = 32'b10010001000101100000001000001011 ^ 32'hf9c75984;
      5'd15: cI7ozekBmfu12 = 32'hf2b3aa10 ^ 32'd2162462033;
      5'd17: cI7ozekBmfu12 = 32'hfba8d4a6 ^ 32'o27634265135 ^ 32'h29f14eee;
      5'd18: cI7ozekBmfu12 = 32'b01001101110110100010101000101001 ^ 32'd2906161017 ^ 32'o35042242373;
      5'd0: cI7ozekBmfu12 = 32'd2427065876 ^ 32'h32dfb430 ^ 32'd2448352559;
      5'b11100: cI7ozekBmfu12 = 32'o20113500275 ^ 32'o23253351161;
      5'b11010: cI7ozekBmfu12 = 32'hd64f63f ^ 32'o33477054234 ^ 32'b10001000000001100111111111000101;
      5'h13: cI7ozekBmfu12 = 32'b11011010001101010010100010001100 ^ 32'b11000101110100010011111001000111 ^ 32'd1101102879;
      5'b00100: cI7ozekBmfu12 = 32'o26774060011 ^ 32'b11010011010010101000000101010011;
      5'o1: cI7ozekBmfu12 = 32'b00111000110101001110010011010010 ^ 32'o3437254022;
      5'b01011: cI7ozekBmfu12 = 32'ha255376d ^ 32'd497586730 ^ 32'b10101100110001001100111011000000;
      5'b01010: cI7ozekBmfu12 = 32'b01100110001001001011101000010010 ^ 32'o11600330143;
      5'o26: cI7ozekBmfu12 = 32'd4006329442 ^ 32'd3621918242;
      5'd16: cI7ozekBmfu12 = 32'b10110101100011011100011101100110 ^ 32'h3b5e545e ^ 32'h9160d6f6;
      5'd3: cI7ozekBmfu12 = 32'd416949840 ^ 32'o10462532570 ^ 32'd1644801955;
      5'd14: cI7ozekBmfu12 = 32'd1290782539 ^ 32'd4086207925 ^ 32'o25520616677;
      5'o24: cI7ozekBmfu12 = 32'd3063480191 ^ 32'd2835015402;
    endcase
  end

  always_ff @(posedge clk_i) begin
    if(zZF) begin
      X5ldx3X4a <= '0;
    end else if (jMTaMbqs055c0zWDyuyX[32'd15091 ^ 32'd28271 ^ 32'o65644 ^ 32'h4036 ^ 32'b00000000000000000110010001100010 ^ 32'o15555]) begin
      X5ldx3X4a <= '0;
    end
    else if(cI7ozekBmfu12[32'o13355 ^ 32'b00000000000000000101111011100001 ^ 32'o44011]) begin
      case(UmLX)
        32'h00: X5ldx3X4a <= data;
        32'h04: X5ldx3X4a <= valid;
        32'h08: X5ldx3X4a <= busy;
        32'h0c: X5ldx3X4a <= baudrate;
        32'h10: X5ldx3X4a <= parity_en;
        32'h14: X5ldx3X4a <= stopbit;
        default: X5ldx3X4a <= X5ldx3X4a;
      endcase
    end
    else begin
      X5ldx3X4a <= X5ldx3X4a;
    end
  end

  always_ff @(posedge clk_i) begin
    if(zZF) begin
      stopbit <= '0;
    end else if (WLGbSSV5YzHmlpmqLI[32'b00000000000000000000010011110011 ^ 32'b00000000000000000111111100110011 ^ 32'h7bc1]) begin
      stopbit <= '0;
    end else if(vBjc8EzRDlz48WXa4k[32'h207b ^ 32'o24252 ^ 32'h7639 ^ 32'h764 ^ 32'o20713 ^ 32'd30353 ^ 32'b00000000000000000010001101000100 ^ 32'o6627]) begin
      stopbit <= FFDK4sD9m7;
    end
    else begin
      stopbit <= stopbit;
    end
  end
  assign q0MK89N8qKhS8mdymRsz = FFDK4sD9m7[0];
  assign pEo = req_i;
endmodule
