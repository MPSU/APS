/* -----------------------------------------------------------------------------
* Project Name   : Architectures of Processor Systems (APS) lab work
* Organization   : National Research University of Electronic Technology (MIET)
* Department     : Institute of Microdevices and Control Systems
* Author(s)      : Andrei Solodovnikov
* Email(s)       : hepoh@org.miet.ru

See https://github.com/MPSU/APS/blob/master/LICENSE file for licensing details.
* ------------------------------------------------------------------------------
*/
module tb_blaster();

  logic          clk_i;
  logic          rst_i;
  logic          rx_i;
  logic          tx_o;
  logic [ 31:0]  instr_addr_o;
  logic [ 31:0]  instr_wdata_o;
  logic          instr_write_enable_o;
  logic [ 31:0]  data_addr_o;
  logic [ 31:0]  data_wdata_o;
  logic          data_write_enable_o;
  logic [ 31:0]  tiff_addr_o;
  logic [127:0]  tiff_wdata_o;
  logic          tiff_write_enable_o;
  logic          core_reset_o;

  logic rx_busy, rx_valid, tx_busy, tx_valid;
  logic [7:0] rx_data, tx_data;

  logic [31:0]   instr_addr_i;
  logic [31:0]   instr_rdata_o;
  logic [31:0]   tiff_addr_i;
  logic [127:0]  tiff_rdata_o;

  logic [3:0] [7:0] flash_addr;
  logic [3:0] [7:0] instr_size;
  logic [3:0] [7:0] instr_size_ack;
  logic [3:0] [7:0] data_size;
  logic [3:0] [7:0] data_size_ack;
  logic [3:0] [7:0] tiff_size;
  logic [3:0] [7:0] tiff_size_ack;

  logic [7:0] instr_mem_byte[$];
  logic [7:0] data_mem_byte[$];
  logic [7:0] tiff_mem_byte [$];

  localparam INIT_MSG_SIZE  = 40;
  localparam MSG_DONE_SIZE  = 57;
  localparam MSG_ACK_SIZE   = 4;

  byte init_str[INIT_MSG_SIZE];
  byte done_str[MSG_DONE_SIZE];

  always #50ns clk_i = !clk_i;

  initial begin
    $timeformat(-9, 2, " ns", 3);
    clk_i = 0;
    rst_i <= 0;
    @(posedge clk_i);
    rst_i <= 1;
    repeat(2) @(posedge clk_i);
    rst_i <= 0;
    instr_size = instr_mem_byte.size();
    data_size  = data_mem_byte.size();
    tiff_size  = tiff_mem_byte.size();
    
/*
    RCV_NEXT_COMMAND
*/
    flash_addr = 32'h0000;
    for(int i = MSG_ACK_SIZE-1; i >= 0; i--) begin
      tx_data = flash_addr[i];
      tx_valid = 1'b1;
      @(posedge clk_i);
      tx_valid = 1'b0;
      @(posedge clk_i);
      while(tx_busy) @(posedge clk_i);
    end

/*
    INIT_MSG
*/
    for(int i = 0; i < INIT_MSG_SIZE; i++) begin
      @(posedge clk_i);
      while(!rx_valid)@(posedge clk_i);
      init_str[i] = rx_data;
    end
    $display("%s", init_str);
    wait(tx_o);
//  ----------------------------------------------

    repeat(10000)@(posedge clk_i);

/*
    RCV_INSTR_SIZE
*/
    for(int i = MSG_ACK_SIZE-1; i >= 0; i--) begin
      tx_data = instr_size[i];
      tx_valid = 1'b1;
      @(posedge clk_i);
      tx_valid = 1'b0;
      @(posedge clk_i);
      while(tx_busy) @(posedge clk_i);
    end
//  ----------------------------------------------


/*
    INSTR_SIZE_ACK
*/
    for(int i = MSG_ACK_SIZE-1; i >= 0; i--) begin
      while(!rx_valid) @(posedge clk_i);
      instr_size_ack[i] = rx_data;
      @(posedge clk_i);
    end
    $display("%h", instr_size);
    assert(instr_size_ack == instr_size)
    else $error("ack: %0h, size: %0h", instr_size_ack, instr_size);
    wait(tx_o);
//  ----------------------------------------------



/*
    INSTR_FLASH
*/
    if(instr_size)repeat(10000)@(posedge clk_i);
    for(int i = instr_size-1; i >=0; i--) begin
      tx_data = instr_mem_byte[i];
      tx_valid = 1'b1;
      @(posedge clk_i);
      tx_valid = 1'b0;
      @(posedge clk_i);
      while(tx_busy) @(posedge clk_i);
    end
//  ----------------------------------------------


/*
    INSTR_FLASH_ACK
*/
    for(int i = 0; i < MSG_DONE_SIZE; i++) begin
      @(posedge clk_i);
      while(!rx_valid)@(posedge clk_i);
      done_str[i] = rx_data;
    end
    $display("%t %s", $time, done_str);
    wait(tx_o);
//  ----------------------------------------------



    repeat(10000)@(posedge clk_i);

/*
    RCV_NEXT_COMMAND
*/  flash_addr = 32'h4000;
    for(int i = MSG_ACK_SIZE-1; i >= 0; i--) begin
      tx_data = flash_addr[i];
      tx_valid = 1'b1;
      @(posedge clk_i);
      tx_valid = 1'b0;
      @(posedge clk_i);
      while(tx_busy) @(posedge clk_i);
    end


/*
    INIT_MSG
*/
    for(int i = 0; i < INIT_MSG_SIZE; i++) begin
      @(posedge clk_i);
      while(!rx_valid)@(posedge clk_i);
      init_str[i] = rx_data;
    end
    $display("%s", init_str);
    wait(tx_o);
//  ----------------------------------------------

/*
    RCV_DATA_SIZE
*/
    for(int i = MSG_ACK_SIZE-1; i >= 0; i--) begin
      tx_data = data_size[i];
      tx_valid = 1'b1;
      @(posedge clk_i);
      tx_valid = 1'b0;
      @(posedge clk_i);
      while(tx_busy) @(posedge clk_i);
    end
//  ----------------------------------------------


/*
    DATA_SIZE_ACK
*/
    for(int i = MSG_ACK_SIZE-1; i >= 0; i--) begin
      while(!rx_valid) @(posedge clk_i);
      data_size_ack[i] = rx_data;
      @(posedge clk_i);
    end
    $display("%h", data_size);
    assert(data_size_ack == data_size)
    else $error("ack: %0h, size: %0h", data_size_ack, data_size);
    wait(tx_o);
//  ----------------------------------------------


/*
    DATA_FLASH
*/
    if(data_size)repeat(10000)@(posedge clk_i);
    for(int i = data_size-1; i >=0; i--) begin
      tx_data = data_mem_byte[i];
      tx_valid = 1'b1;
      @(posedge clk_i);
      tx_valid = 1'b0;
      @(posedge clk_i);
      while(tx_busy) @(posedge clk_i);
    end
//  ----------------------------------------------


/*
    DATA_FLASH_ACK
*/
    for(int i = 0; i < MSG_DONE_SIZE; i++) begin
      @(posedge clk_i);
      while(!rx_valid)@(posedge clk_i);
      done_str[i] = rx_data;
    end
    $display("%t %s", $time, done_str);
    wait(tx_o);
//  ----------------------------------------------
    repeat(10000)@(posedge clk_i);


/*
    RCV_NEXT_COMMAND
*/  flash_addr = 32'h0800_0000;
    for(int i = MSG_ACK_SIZE-1; i >= 0; i--) begin
      tx_data = flash_addr[i];
      tx_valid = 1'b1;
      @(posedge clk_i);
      tx_valid = 1'b0;
      @(posedge clk_i);
      while(tx_busy) @(posedge clk_i);
    end

/*
    INIT_MSG
*/
    for(int i = 0; i < INIT_MSG_SIZE; i++) begin
      @(posedge clk_i);
      while(!rx_valid)@(posedge clk_i);
      init_str[i] = rx_data;
    end
    $display("%s", init_str);
    wait(tx_o);
//  ----------------------------------------------

/*
    RCV_TIFF_SIZE
*/
    for(int i = MSG_ACK_SIZE-1; i >= 0; i--) begin
      tx_data = tiff_size[i];
      tx_valid = 1'b1;
      @(posedge clk_i);
      tx_valid = 1'b0;
      @(posedge clk_i);
      while(tx_busy) @(posedge clk_i);
    end
//  ----------------------------------------------


/*
    TIFF_SIZE_ACK
*/
    for(int i = MSG_ACK_SIZE-1; i >= 0; i--) begin
      while(!rx_valid) @(posedge clk_i);
      tiff_size_ack[i] = rx_data;
      @(posedge clk_i);
    end
    $display("%h", tiff_size);
    assert(tiff_size_ack == tiff_size)
    else $display("ack: %0h, size: %0h", tiff_size_ack, tiff_size);
    wait(tx_o);
//  ----------------------------------------------



/*
    TIFF_FLASH
*/
    if(tiff_size)repeat(10000)@(posedge clk_i);
    for(int i = tiff_size-1; i >=0; i--) begin
      tx_data = tiff_mem_byte[i];
      tx_valid = 1'b1;
      @(posedge clk_i);
      tx_valid = 1'b0;
      @(posedge clk_i);
      while(tx_busy) @(posedge clk_i);
    end
//  ----------------------------------------------


/*
    TIFF_FLASH_ACK, FINISH
*/
    for(int i = 0; i < MSG_DONE_SIZE; i++) begin
      @(posedge clk_i);
      while(!rx_valid)@(posedge clk_i);
      done_str[i] = rx_data;
    end
    $display("%t %s", $time, done_str);
    wait(!rx_busy)
    @(posedge clk_i)

/*
    RCV_NEXT_COMMAND
*/  flash_addr = 32'hFFFF_FFFF;
    for(int i = MSG_ACK_SIZE-1; i >= 0; i--) begin
      tx_data = flash_addr[i];
      tx_valid = 1'b1;
      @(posedge clk_i);
      tx_valid = 1'b0;
      @(posedge clk_i);
      while(tx_busy) @(posedge clk_i);
    end

    assert(!core_reset_o)
    else $error("reset is not equal zero at the end");
//  ----------------------------------------------

    repeat(10000)@(posedge clk_i);

    $finish();
  end


  bluster blust(.*);

  uart_rx rx(
  .clk_i      (clk_i      ),
  .rst_i      (rst_i      ),
  .rx_i       (tx_o       ),
  .busy_o     (rx_busy    ),
  .baudrate_i (17'd115200 ),
  .parity_en_i(1'b1       ),
  .stopbit_i  (1'b1       ),
  .rx_data_o  (rx_data    ),
  .rx_valid_o (rx_valid   )
);

uart_tx tx(
  .clk_i      (clk_i      ),
  .rst_i      (rst_i      ),
  .tx_o       (rx_i       ),
  .busy_o     (tx_busy    ),
  .baudrate_i (17'd115200 ),
  .parity_en_i(1'b1       ),
  .stopbit_i  (1'b1       ),
  .tx_data_i  (tx_data    ),
  .tx_valid_i (tx_valid   )
);

  rw_instr_mem imem(
    .clk_i         (clk_i               ) ,
    .read_addr_i   (instr_addr_i        ) ,
    .read_data_o   (instr_rdata_o       ) ,
    .write_addr_i  (instr_addr_o        ) ,
    .write_data_i  (instr_wdata_o       ) ,
    .write_enable_i(instr_write_enable_o)
  );

  ext_mem dmem(
    .clk_i          (clk_i              ),
    .mem_req_i      (data_addr_o[31:24] == 0),
    .write_enable_i (data_write_enable_o),
    .byte_enable_i  (4'b1111            ),
    .addr_i         (data_addr_o        ),
    .write_data_i   (data_wdata_o       ),
    .read_data_o    (),
    .ready_o        ()
  );

  ext_mem tmem(
    .clk_i          (clk_i              ),
    .mem_req_i      (data_addr_o[31:24] == 8),
    .write_enable_i (data_write_enable_o),
    .byte_enable_i  (4'b1111            ),
    .addr_i         (data_addr_o        ),
    .write_data_i   (data_wdata_o       ),
    .read_data_o    (),
    .ready_o        ()
  );

initial instr_mem_byte = {
8'h93, 8'h00, 8'h10, 8'h00, 8'h37, 8'h01, 8'h00, 8'h06, 8'hB7, 8'hC1, 8'h01, 8'h00, 8'h93, 8'h81, 8'h01, 8'h20,
8'h23, 8'h26, 8'h31, 8'h00, 8'h13, 8'h02, 8'h10, 8'h00, 8'h23, 8'h28, 8'h41, 8'h00, 8'h93, 8'h02, 8'h10, 8'h00,
8'h93, 8'h80, 8'h10, 8'h00, 8'h83, 8'h23, 8'h81, 8'h00, 8'h63, 8'h14, 8'h70, 8'h00, 8'h6F, 8'h00, 8'h00, 8'h00,
8'h6F, 8'h00, 8'h00, 8'h00, 8'h23, 8'h20, 8'h11, 8'h00, 8'h6F, 8'h00, 8'h00, 8'h00
};

initial #1 data_mem_byte = instr_mem_byte;

initial tiff_mem_byte = {
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000101, 8'b00000101, 8'b00000101, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00010010, 8'b00010010, 8'b00111111, 8'b00010010, 8'b00010010, 8'b00010010, 8'b00111111, 8'b00010010, 8'b00010010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000100, 8'b00001110, 8'b00010001, 8'b00010001, 8'b00000001, 8'b00001110, 8'b00010000, 8'b00010000, 8'b00010001, 8'b00010001, 8'b00001110, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000010, 8'b00000101, 8'b01000101, 8'b00100010, 8'b00010000, 8'b00001000, 8'b00000100, 8'b00100010, 8'b01010001, 8'b01010000, 8'b00100000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00001100, 8'b00010010, 8'b00010010, 8'b00010010, 8'b01001100, 8'b01001010, 8'b00110001, 8'b00100001, 8'b00110001, 8'b01001110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00010010, 8'b00001100, 8'b00111111, 8'b00001100, 8'b00010010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000100, 8'b00011111, 8'b00000100, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00010000, 8'b00010000, 8'b00001000, 8'b00001000, 8'b00000100, 8'b00000100, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00110001, 8'b00101001, 8'b00101001, 8'b00100101, 8'b00100101, 8'b00100011, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00001000, 8'b00001100, 8'b00001010, 8'b00001001, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100000, 8'b00010000, 8'b00001000, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100000, 8'b00100000, 8'b00011100, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00010000, 8'b00011000, 8'b00010100, 8'b00010010, 8'b00010001, 8'b00111111, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00111111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00011111, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011100, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00111111, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00010000, 8'b00001000, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00111110, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00010000, 8'b00001000, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00000010, 8'b00000100, 8'b00001000, 8'b00010000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b00000000, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000100, 8'b00001000, 8'b00010000, 8'b00001000, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100000, 8'b00010000, 8'b00001000, 8'b00000100, 8'b00000000, 8'b00000100, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b01000010, 8'b10011001, 8'b10100001, 8'b10111001, 8'b10100101, 8'b01111001, 8'b00000010, 8'b01111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00111111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00001111, 8'b00010001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00010001, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00111111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00001111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00111111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00001111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00111001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00111111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00100001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00100001, 8'b00100001, 8'b00010001, 8'b00001001, 8'b00000111, 8'b00001001, 8'b00010001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b01000001, 8'b01100011, 8'b01010101, 8'b01001001, 8'b01001001, 8'b01000001, 8'b01000001, 8'b01000001, 8'b01000001, 8'b01000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00100001, 8'b00100011, 8'b00100101, 8'b00101001, 8'b00110001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00101001, 8'b00110001, 8'b00111110, 8'b00100000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011111, 8'b00010001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00000001, 8'b00000010, 8'b00001100, 8'b00010000, 8'b00100000, 8'b00100000, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b01111111, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b01000001, 8'b01000001, 8'b01000001, 8'b01000001, 8'b00100010, 8'b00100010, 8'b00010100, 8'b00010100, 8'b00001000, 8'b00001000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b01000001, 8'b01000001, 8'b01000001, 8'b01000001, 8'b01001001, 8'b01001001, 8'b01001001, 8'b01010101, 8'b01100011, 8'b01000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00010010, 8'b00001100, 8'b00001100, 8'b00010010, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b01000001, 8'b01000001, 8'b00100010, 8'b00100010, 8'b00010100, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00111111, 8'b00100000, 8'b00100000, 8'b00010000, 8'b00001000, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000100, 8'b00000100, 8'b00001000, 8'b00001000, 8'b00010000, 8'b00010000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000111, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000100, 8'b00001010, 8'b00010001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00100000, 8'b00111110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00111110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00111110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00111110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00111111, 8'b00000001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011100, 8'b00100010, 8'b00000010, 8'b00000010, 8'b00001111, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00110001, 8'b00101110, 8'b00100000, 8'b00100001, 8'b00011110, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00010000, 8'b00000000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010001, 8'b00010001, 8'b00001110, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00100001, 8'b00100001, 8'b00010001, 8'b00001111, 8'b00010001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00110111, 8'b01001001, 8'b01001001, 8'b01001001, 8'b01001001, 8'b01001001, 8'b01000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00111110, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011101, 8'b00000011, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00000001, 8'b00011110, 8'b00100000, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000100, 8'b00011111, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00011000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00111110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000001, 8'b01000001, 8'b00100010, 8'b00100010, 8'b00010100, 8'b00010100, 8'b00001000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000001, 8'b01000001, 8'b01001001, 8'b01001001, 8'b01001001, 8'b01010101, 8'b00100010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000001, 8'b00100010, 8'b00010100, 8'b00001000, 8'b00010100, 8'b00100010, 8'b01000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00110001, 8'b00101110, 8'b00100000, 8'b00010000, 8'b00001111, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b00010000, 8'b00001000, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011000, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000011, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00011000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000011, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00011000, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000011, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00100110, 8'b00011001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000011, 8'b00000101, 8'b00000101, 8'b00000011, 8'b00000000, 8'b00001100, 8'b00001100, 8'b00000100, 8'b00101100, 8'b00100000, 8'b00100000, 8'b01100000, 8'b00000000, 8'b00000000, 8'b00000000
};

endmodule


module rw_tiff_mem(
  input  logic         clk_i,
  input  logic [ 31:0] addr_i,
  output logic [127:0] read_data_o,

  input  logic [ 31:0] write_addr_i,
  input  logic [127:0] write_data_i,
  input  logic         write_enable_i
);

logic [127:0] rom [256];

assign read_data_o = rom[addr_i];

always_ff @(posedge clk_i) begin
  if(write_enable_i) begin
    rom[write_addr_i] <= write_data_i;
  end
end

endmodule