/* -----------------------------------------------------------------------------
* Project Name   : Architectures of Processor Systems (APS) lab work
* Organization   : National Research University of Electronic Technology (MIET)
* Department     : Institute of Microdevices and Control Systems
* Author(s)      : Andrei Solodovnikov
* Email(s)       : hepoh@org.miet.ru

See https://github.com/MPSU/APS/blob/master/LICENSE file for licensing details.
* ------------------------------------------------------------------------------
*/
module tb_top_asic();

  logic        clk10mhz_i;
  logic        aresetn_i;
  logic        rx_i;
  logic        tx_o;
  logic          clk_i;
  logic          rst_i;

  assign aresetn_i = !rst_i;
  assign clk10mhz_i = clk_i;

  logic rx_busy, rx_valid, tx_busy, tx_valid;
  logic [7:0] rx_data, tx_data;

  logic [3:0] [7:0] instr_size_ack;
  logic [3:0] [7:0] data_size_ack;
  logic [3:0] [7:0] tiff_size = 32'd0;
  logic [3:0] [7:0] tiff_size_ack;
  byte init_str[6];
  byte done_str[10];
  logic [7:0] instr_mem_byte[];
  logic [7:0] data_mem_byte[];
  logic [3:0] [7:0] instr_size;
  logic [3:0] [7:0] data_size;

  initial begin
    // $readmemh("tb_coremark_instr.mem", instr_mem_byte);
    // $readmemh("tb_coremark_data.mem", data_mem_byte);
    // instr_size = instr_mem_byte.size();
    // data_size  = data_mem_byte.size();
    instr_size = 0;
    data_size  = 0;
  end

  logic [7:0] tiff_mem_byte [2048];

  localparam INIT_MSG_SIZE  = 6;
  localparam MSG_DONE_SIZE  = 10;
  localparam MSG_ACK_SIZE   = 4;

  always #50ns clk_i = !clk_i;

  byte coremark_msg[103];
  integer coremark_cntr;

  initial begin
    $timeformat(-9, 2, " ns", 3);
    clk_i = 0;
    rst_i <= 0;
    @(posedge clk_i);
    rst_i <= 1;
    repeat(2) @(posedge clk_i);
    rst_i <= 0;

/*
    INIT_MSG
*/
    for(int i = 0; i < INIT_MSG_SIZE; i++) begin
      @(posedge clk_i);
      while(!rx_valid)@(posedge clk_i);
      init_str[i] = rx_data;
    end
    $display("%s", init_str);
    wait(tx_o);
//  ----------------------------------------------

    repeat(10000)@(posedge clk_i);

/*
    IDLE, RCV_INSTR_SIZE
*/
    for(int i = MSG_ACK_SIZE-1; i >= 0; i--) begin
      tx_data = instr_size[i];
      tx_valid = 1'b1;
      @(posedge clk_i);
      tx_valid = 1'b0;
      @(posedge clk_i);
      while(tx_busy) @(posedge clk_i);
    end
//  ----------------------------------------------


/*
    INSTR_SIZE_ACK
*/
    for(int i = MSG_ACK_SIZE-1; i >= 0; i--) begin
      while(!rx_valid) @(posedge clk_i);
      instr_size_ack[i] = rx_data;
      @(posedge clk_i);
    end
    assert(instr_size_ack == instr_size)
    else $error("ack: %0h, size: %0h", instr_size_ack, instr_size);
    wait(tx_o);
//  ----------------------------------------------



/*
    INSTR_FLASH
*/
    if(instr_size)repeat(10000)@(posedge clk_i);
    for(int i = instr_size-1; i >=0; i--) begin
      tx_data = instr_mem_byte[i];
      tx_valid = 1'b1;
      @(posedge clk_i);
      tx_valid = 1'b0;
      @(posedge clk_i);
      while(tx_busy) @(posedge clk_i);
    end
//  ----------------------------------------------


/*
    INSTR_FLASH_ACK
*/
    for(int i = 0; i < MSG_DONE_SIZE; i++) begin
      @(posedge clk_i);
      while(!rx_valid)@(posedge clk_i);
      done_str[i] = rx_data;
    end
    $display("%t %s", $time, done_str);
    wait(tx_o);
//  ----------------------------------------------



    repeat(10000)@(posedge clk_i);



/*
    RCV_DATA_SIZE
*/
    for(int i = MSG_ACK_SIZE-1; i >= 0; i--) begin
      tx_data = data_size[i];
      tx_valid = 1'b1;
      @(posedge clk_i);
      tx_valid = 1'b0;
      @(posedge clk_i);
      while(tx_busy) @(posedge clk_i);
    end
//  ----------------------------------------------


/*
    DATA_SIZE_ACK
*/
    for(int i = MSG_ACK_SIZE-1; i >= 0; i--) begin
      while(!rx_valid) @(posedge clk_i);
      data_size_ack[i] = rx_data;
      @(posedge clk_i);
    end
    assert(data_size_ack == data_size)
    else $error("ack: %0h, size: %0h", data_size_ack, data_size);
    wait(tx_o);
//  ----------------------------------------------


/*
    DATA_FLASH
*/
    if(data_size)repeat(10000)@(posedge clk_i);
    for(int i = data_size-1; i >=0; i--) begin
      tx_data = data_mem_byte[i];
      tx_valid = 1'b1;
      @(posedge clk_i);
      tx_valid = 1'b0;
      @(posedge clk_i);
      while(tx_busy) @(posedge clk_i);
    end
//  ----------------------------------------------


/*
    DATA_FLASH_ACK
*/
    for(int i = 0; i < MSG_DONE_SIZE; i++) begin
      @(posedge clk_i);
      while(!rx_valid)@(posedge clk_i);
      done_str[i] = rx_data;
    end
    $display("%t %s", $time, done_str);
    wait(tx_o);
//  ----------------------------------------------
    repeat(10000)@(posedge clk_i);





/*
    RCV_TIFF_SIZE
*/
    for(int i = MSG_ACK_SIZE-1; i >= 0; i--) begin
      tx_data = tiff_size[i];
      tx_valid = 1'b1;
      @(posedge clk_i);
      tx_valid = 1'b0;
      @(posedge clk_i);
      while(tx_busy) @(posedge clk_i);
    end
//  ----------------------------------------------


/*
    TIFF_SIZE_ACK
*/
    for(int i = MSG_ACK_SIZE-1; i >= 0; i--) begin
      while(!rx_valid) @(posedge clk_i);
      tiff_size_ack[i] = rx_data;
      @(posedge clk_i);
    end
    assert(tiff_size_ack == tiff_size)
    else $display("ack: %0h, size: %0h", tiff_size_ack, tiff_size);
    wait(tx_o);
//  ----------------------------------------------



/*
    TIFF_FLASH
*/
    if(tiff_size)repeat(10000)@(posedge clk_i);
    for(int i = tiff_size-1; i >=0; i--) begin
      tx_data = tiff_mem_byte[i];
      tx_valid = 1'b1;
      @(posedge clk_i);
      tx_valid = 1'b0;
      @(posedge clk_i);
      while(tx_busy) @(posedge clk_i);
    end
//  ----------------------------------------------


/*
    TIFF_FLASH_ACK, FINISH
*/
    for(int i = 0; i < MSG_DONE_SIZE; i++) begin
      @(posedge clk_i);
      while(!rx_valid)@(posedge clk_i);
      done_str[i] = rx_data;
    end
    $display("%t %s", $time, done_str);
    wait(!rx_busy)
    @(posedge clk_i)
    // assert(!pc_stall_o)
    // else $error("stall is not equal zero at the end");
//  ----------------------------------------------

    repeat(10000)@(posedge clk_i);
    coremark_cntr = 0;
    coremark_msg = {32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32};
    forever begin
      @(posedge clk_i);
      if(rx_valid) begin
        if((rx_data == 10) | (rx_data == 13)) begin
          $display("%s", coremark_msg);
          coremark_cntr = 0;
          coremark_msg = {32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32};
        end
        else begin
          coremark_msg[coremark_cntr] = rx_data;
          coremark_cntr++;
        end
      end
    end
    // $finish();
  end


  riscv_top_asic DUT(.clk10mhz_i, .aresetn_i, .rx_i, .tx_o);

  uart_rx rx(
  .clk_i      (clk_i      ),
  .rst_i      (rst_i      ),
  .rx_i       (tx_o       ),
  .busy_o     (rx_busy    ),
  .baudrate_i (17'd115200 ),
  .parity_en_i(1'b1       ),
  .stopbit_i  (1'b1       ),
  .rx_data_o  (rx_data    ),
  .rx_valid_o (rx_valid   )
);

uart_tx tx(
  .clk_i      (clk_i      ),
  .rst_i      (rst_i      ),
  .tx_o       (rx_i       ),
  .busy_o     (tx_busy    ),
  .baudrate_i (17'd115200 ),
  .parity_en_i(1'b1       ),
  .stopbit_i  (1'b1       ),
  .tx_data_i  (tx_data    ),
  .tx_valid_i (tx_valid   )
);


initial tiff_mem_byte = {
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00011110,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000101, 8'b00000101, 8'b00000101, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00010010, 8'b00010010, 8'b00111111, 8'b00010010, 8'b00010010, 8'b00010010, 8'b00111111, 8'b00010010, 8'b00010010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000100, 8'b00001110, 8'b00010001, 8'b00010001, 8'b00000001, 8'b00001110, 8'b00010000, 8'b00010000, 8'b00010001, 8'b00010001, 8'b00001110, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000010, 8'b00000101, 8'b01000101, 8'b00100010, 8'b00010000, 8'b00001000, 8'b00000100, 8'b00100010, 8'b01010001, 8'b01010000, 8'b00100000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00001100, 8'b00010010, 8'b00010010, 8'b00010010, 8'b01001100, 8'b01001010, 8'b00110001, 8'b00100001, 8'b00110001, 8'b01001110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00010010, 8'b00001100, 8'b00111111, 8'b00001100, 8'b00010010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000100, 8'b00011111, 8'b00000100, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00010000, 8'b00010000, 8'b00001000, 8'b00001000, 8'b00000100, 8'b00000100, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00110001, 8'b00101001, 8'b00101001, 8'b00100101, 8'b00100101, 8'b00100011, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00001000, 8'b00001100, 8'b00001010, 8'b00001001, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100000, 8'b00010000, 8'b00001000, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100000, 8'b00100000, 8'b00011100, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00010000, 8'b00011000, 8'b00010100, 8'b00010010, 8'b00010001, 8'b00111111, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00111111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00011111, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011100, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00111111, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00010000, 8'b00001000, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00111110, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000010, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00010000, 8'b00001000, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00000010, 8'b00000100, 8'b00001000, 8'b00010000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b00000000, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000010, 8'b00000100, 8'b00001000, 8'b00010000, 8'b00001000, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100000, 8'b00010000, 8'b00001000, 8'b00000100, 8'b00000000, 8'b00000100, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b01000010, 8'b10011001, 8'b10100001, 8'b10111001, 8'b10100101, 8'b01111001, 8'b00000010, 8'b01111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00111111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00001111, 8'b00010001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00010001, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00111111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00001111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00111111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00001111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00111001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00111111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00100001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00100001, 8'b00100001, 8'b00010001, 8'b00001001, 8'b00000111, 8'b00001001, 8'b00010001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b01000001, 8'b01100011, 8'b01010101, 8'b01001001, 8'b01001001, 8'b01000001, 8'b01000001, 8'b01000001, 8'b01000001, 8'b01000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00100001, 8'b00100011, 8'b00100101, 8'b00101001, 8'b00110001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00101001, 8'b00110001, 8'b00111110, 8'b00100000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011111, 8'b00010001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00000001, 8'b00000010, 8'b00001100, 8'b00010000, 8'b00100000, 8'b00100000, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b01111111, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b01000001, 8'b01000001, 8'b01000001, 8'b01000001, 8'b00100010, 8'b00100010, 8'b00010100, 8'b00010100, 8'b00001000, 8'b00001000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b01000001, 8'b01000001, 8'b01000001, 8'b01000001, 8'b01001001, 8'b01001001, 8'b01001001, 8'b01010101, 8'b01100011, 8'b01000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00010010, 8'b00001100, 8'b00001100, 8'b00010010, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b01000001, 8'b01000001, 8'b00100010, 8'b00100010, 8'b00010100, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00001000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00111111, 8'b00100000, 8'b00100000, 8'b00010000, 8'b00001000, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00000001, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000010, 8'b00000100, 8'b00000100, 8'b00001000, 8'b00001000, 8'b00010000, 8'b00010000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000111, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000100, 8'b00001010, 8'b00010001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00100000, 8'b00111110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00111110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00111110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00111110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00111111, 8'b00000001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011100, 8'b00100010, 8'b00000010, 8'b00000010, 8'b00001111, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00110001, 8'b00101110, 8'b00100000, 8'b00100001, 8'b00011110, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00010000, 8'b00000000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010000, 8'b00010001, 8'b00010001, 8'b00001110, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00100001, 8'b00100001, 8'b00010001, 8'b00001111, 8'b00010001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00110111, 8'b01001001, 8'b01001001, 8'b01001001, 8'b01001001, 8'b01001001, 8'b01000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011111, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00011111, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111110, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00111110, 8'b00100000, 8'b00100000, 8'b00100000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011101, 8'b00000011, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00100001, 8'b00000001, 8'b00011110, 8'b00100000, 8'b00100001, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000100, 8'b00000100, 8'b00011111, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00011000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00111110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000001, 8'b01000001, 8'b00100010, 8'b00100010, 8'b00010100, 8'b00010100, 8'b00001000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000001, 8'b01000001, 8'b01001001, 8'b01001001, 8'b01001001, 8'b01010101, 8'b00100010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000001, 8'b00100010, 8'b00010100, 8'b00001000, 8'b00010100, 8'b00100010, 8'b01000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00100001, 8'b00110001, 8'b00101110, 8'b00100000, 8'b00010000, 8'b00001111, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b00010000, 8'b00001000, 8'b00000100, 8'b00000010, 8'b00000001, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00011000, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000011, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00011000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00000011, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00011000, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000100, 8'b00000011, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000000, 8'b00100110, 8'b00011001, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
8'b00000000, 8'b00000011, 8'b00000101, 8'b00000101, 8'b00000011, 8'b00000000, 8'b00001100, 8'b00001100, 8'b00000100, 8'b00101100, 8'b00100000, 8'b00100000, 8'b01100000, 8'b00000000, 8'b00000000, 8'b00000000
};

endmodule


module rw_tiff_mem(
  input  logic         clk_i,
  input  logic [ 31:0] addr_i,
  output logic [127:0] read_data_o,

  input  logic [ 31:0] write_addr_i,
  input  logic [127:0] write_data_i,
  input  logic         write_enable_i
);

logic [127:0] rom [256];

assign read_data_o = rom[addr_i];

always_ff @(posedge clk_i) begin
  if(write_enable_i) begin
    rom[write_addr_i] <= write_data_i;
  end
end

endmodule