module uart_tx_sb_ctrl(
/*
    Часть интерфейса модуля, отвечающая за подключение к системной шине
*/
  input  logic          clk_i,
  input  logic          rst_i,
  input  logic [31:0]   addr_i,
  input  logic          req_i,
  input  logic [31:0]   write_data_i,
  input  logic          write_enable_i,
  output logic [31:0]   read_data_o,

/*
    Часть интерфейса модуля, отвечающая за подключение передающему,
    входные данные по UART
*/
  output logic          tx_o
);

  logic [31:0]   Y2pd;
  assign Y2pd = addr_i;
  logic          Uzd;
  assign Uzd = req_i;
  logic [31:0]   ra2VgcBEzc;
  assign ra2VgcBEzc = write_data_i;
  logic          Gdxya89mlifb;
  assign Gdxya89mlifb = write_enable_i;
  logic [31:0]   eCNnNC8kn;
  assign read_data_o = eCNnNC8kn;

  logic [16:0] baudrate;
  logic parity_en;
  logic [1:0] stopbit;
  logic [7:0] data;
  logic lQ5IWH22X, busy;
  logic cWdgq;

  logic [31:0] gUruyn1hzjChHha47v;

  logic CCdflm;

  logic YAhtnxC5bxEVGCn;

  logic B4zEGLaAwyO6;
  assign B4zEGLaAwyO6 = (ra2VgcBEzc == (32'd4078277091 ^ 32'b10101100000110001101001101010101 ^ 32'b01011111000011010100001010110111));

  assign cWdgq = lQ5IWH22X && CCdflm;

  always_comb begin
    case ({YAhtnxC5bxEVGCn, parity_en, B4zEGLaAwyO6, Gdxya89mlifb, cWdgq, Uzd})
      6'o64: gUruyn1hzjChHha47v = 32'o3402527443 ^ 32'hcdb0b047 ^ 32'b11100110100100001110110111001111;
      6'b100001: gUruyn1hzjChHha47v = 32'o27066366252 ^ 32'h8ff31e01;
      6'd38: gUruyn1hzjChHha47v = 32'he725369b ^ 32'd3490694192;
      6'o51: gUruyn1hzjChHha47v = 32'b10100100100101000011100000010101 ^ 32'd873175144 ^ 32'ha7b552d6;
      6'd11: gUruyn1hzjChHha47v = 32'o20141437101 ^ 32'b01110010101100000001010111001011 ^ 32'hc41cd921;
      6'd7: gUruyn1hzjChHha47v = 32'hddbe52f8 ^ 32'o27325210576 ^ 32'o12160330455;
      6'd13: gUruyn1hzjChHha47v = 32'd1669352754 ^ 32'b10010000101000010110011100010001 ^ 32'o30402754210;
      6'h35: gUruyn1hzjChHha47v = 32'd753523049 ^ 32'o3360625702;
      6'h1d: gUruyn1hzjChHha47v = 32'd2485651753 ^ 32'h42d40d00 ^ 32'he1d6f682;
      6'b000000: gUruyn1hzjChHha47v = 32'ha78b18c4 ^ 32'h90a1ea6f;
      6'h15: gUruyn1hzjChHha47v = 32'hd2369660 ^ 32'd2572713286 ^ 32'd2084837773;
      6'd12: gUruyn1hzjChHha47v = 32'o5577654627 ^ 32'h1ad5ab3c;
      6'b101101: gUruyn1hzjChHha47v = 32'b00010000100110110101101001010011 ^ 32'b11111010100001011100000010011010 ^ 32'o33515064146;
      6'b000110: gUruyn1hzjChHha47v = 32'd1040857706 ^ 32'o1110144301;
      6'b011011: gUruyn1hzjChHha47v = 32'b10110111110110100100110000101000 ^ 32'o20074137203;
      6'b110010: gUruyn1hzjChHha47v = 32'b01011110110010010001000000110000 ^ 32'd487764676 ^ 32'h74f1505f;
      6'h8: gUruyn1hzjChHha47v = 32'b10110010011001110110001101001011 ^ 32'h2db361a5 ^ 32'ha8fef045;
      6'b000101: gUruyn1hzjChHha47v = 32'o31503752604 ^ 32'o10106767035 ^ 32'o27317544462;
      6'd61: gUruyn1hzjChHha47v = 32'h6ef7de81 ^ 32'd3655107485 ^ 32'o20000327663;
      6'd2: gUruyn1hzjChHha47v = 32'b01010110010011101001010010111010 ^ 32'd2088043796 ^ 32'b00011101000100010110001100000101;
      6'b111001: gUruyn1hzjChHha47v = 32'b00001110010001101000111101110111 ^ 32'b00111001011011000111110111011100;
      6'b101010: gUruyn1hzjChHha47v = 32'o25173424252 ^ 32'o34740512255 ^ 32'b01111001010001100100111010101100;
      6'b111111: gUruyn1hzjChHha47v = 32'h5739120f ^ 32'b01100000000100111110000010100000;
      6'd3: gUruyn1hzjChHha47v = 32'o10473305327 ^ 32'o30333052103 ^ 32'b10110000101010110010110000111111;
      6'd25: gUruyn1hzjChHha47v = 32'o11154673764 ^ 32'b01011100111111001101010101001001 ^ 32'd577064982;
      6'd62: gUruyn1hzjChHha47v = 32'o22113121447 ^ 32'ha606518c;
      6'o61: gUruyn1hzjChHha47v = 32'o7375044016 ^ 32'b10110110111110100011011101010011 ^ 32'b10111010001001001000110111110110;
      6'b100010: gUruyn1hzjChHha47v = 32'hfbae602c ^ 32'o33656154567 ^ 32'b00010010001111000100101111110000;
      6'b011110: gUruyn1hzjChHha47v = 32'h2d745bbe ^ 32'h1a5ea915;
      6'h2c: gUruyn1hzjChHha47v = 32'o4304655270 ^ 32'h1439a813;
      6'b010000: gUruyn1hzjChHha47v = 32'h202a19d6 ^ 32'h1700eb7d;
      6'h38: gUruyn1hzjChHha47v = 32'b00101001000100110000110101111001 ^ 32'd2139263367 ^ 32'o14156667125;
      6'o72: gUruyn1hzjChHha47v = 32'h8a37e93 ^ 32'o7742306070;
      6'd26: gUruyn1hzjChHha47v = 32'o17207557126 ^ 32'he574e1c1 ^ 32'ha840cd3c;
      6'd39: gUruyn1hzjChHha47v = 32'hec113b20 ^ 32'd3678128523;
      6'o4: gUruyn1hzjChHha47v = 32'b00000011000010100000100111010000 ^ 32'd874576763;
      6'o57: gUruyn1hzjChHha47v = 32'h5fae971f ^ 32'd4027033477 ^ 32'b10011000100000111100001000110101;
      6'b010111: gUruyn1hzjChHha47v = 32'hc68c2bb2 ^ 32'o13116704315 ^ 32'd2828882388;
      6'b001010: gUruyn1hzjChHha47v = 32'b11101001111011100010001111110010 ^ 32'o33661150531;
      6'b100101: gUruyn1hzjChHha47v = 32'd476563992 ^ 32'b00101011010011010011100010110011;
      6'b101011: gUruyn1hzjChHha47v = 32'h656e2f0f ^ 32'o3171371546 ^ 32'o11350227302;
      6'o73: gUruyn1hzjChHha47v = 32'hdf65c32d ^ 32'b11011000001001010011110011000111 ^ 32'b00110000011010100000110101000001;
      6'b100100: gUruyn1hzjChHha47v = 32'o4613212043 ^ 32'b00010001000001111110011010001000;
      6'h28: gUruyn1hzjChHha47v = 32'b00001111011110110111101101101111 ^ 32'b01111001011110011000010110011110 ^ 32'o10112006132;
      6'o22: gUruyn1hzjChHha47v = 32'o30661233146 ^ 32'd4059022541;
      6'o56: gUruyn1hzjChHha47v = 32'b10010010110111111110110011101111 ^ 32'd1889097106 ^ 32'o32533045726;
      6'b010110: gUruyn1hzjChHha47v = 32'hae0ac991 ^ 32'b11111101110100010001101100110001 ^ 32'h64f1200b;
      6'b000001: gUruyn1hzjChHha47v = 32'd3557726626 ^ 32'd3810814729;
      6'o30: gUruyn1hzjChHha47v = 32'he3e64780 ^ 32'o1365375222 ^ 32'hdf194fb9;
      6'h1c: gUruyn1hzjChHha47v = 32'd2543563122 ^ 32'ha0b143d9;
      6'b110111: gUruyn1hzjChHha47v = 32'ha18a7aa4 ^ 32'b11010101001111100000100111100110 ^ 32'b01000011100111101000000111101001;
      6'b111100: gUruyn1hzjChHha47v = 32'o23306143705 ^ 32'd1638481191 ^ 32'hcd9b0849;
      6'd17: gUruyn1hzjChHha47v = 32'd3809328172 ^ 32'o23771224041 ^ 32'o11360463246;
      6'b110011: gUruyn1hzjChHha47v = 32'b11111110101100011011010001001100 ^ 32'b11001001100110110100011011100111;
      6'o40: gUruyn1hzjChHha47v = 32'd3206040973 ^ 32'hee2f1184 ^ 32'd1713221282;
      6'h14: gUruyn1hzjChHha47v = 32'd309581887 ^ 32'o2520203713 ^ 32'o6006026537;
      6'h1f: gUruyn1hzjChHha47v = 32'o17336311417 ^ 32'o36547100451 ^ 32'd3117408397;
      6'b001111: gUruyn1hzjChHha47v = 32'o20563214357 ^ 32'h4e49558a ^ 32'b11111100101011101011111111001110;
      6'b110000: gUruyn1hzjChHha47v = 32'h7f8d3900 ^ 32'h48a7cbab;
      6'o23: gUruyn1hzjChHha47v = 32'h3816ce0f ^ 32'h80dd164 ^ 32'b00000111001100011110110111000000;
      6'b110110: gUruyn1hzjChHha47v = 32'd3703086281 ^ 32'o35344467142;
      6'o16: gUruyn1hzjChHha47v = 32'b10010110111001010000011110011110 ^ 32'b10100001110011111111010100110101;
      6'b001001: gUruyn1hzjChHha47v = 32'h76796130 ^ 32'd3942942889 ^ 32'b10101010010101110001101100110010;
      6'o43: gUruyn1hzjChHha47v = 32'd1699059059 ^ 32'o12233663730;

      default: gUruyn1hzjChHha47v = 32'hdead_dead;
    endcase
  end
  assign lQ5IWH22X  = Uzd &  Gdxya89mlifb;
  uart_tx tx(
    .clk_i      (clk_i),
    .rst_i      (rst_i),
    .tx_o       (tx_o),
    .busy_o     (busy),
    .baudrate_i (baudrate),
    .parity_en_i(parity_en),
    .stopbit_i  (stopbit),
    .tx_data_i  (ra2VgcBEzc[7:0]),
    .tx_valid_i (cWdgq)
  );
  logic [31:0] j22I6zJCUqZP;
  assign YAhtnxC5bxEVGCn = (Y2pd == (32'd2261272313 ^ 32'd4194190281 ^ 32'o17715402424));

  logic [31:0] Mmiaej2;
  always_comb begin
    case ({YAhtnxC5bxEVGCn, parity_en, busy, Gdxya89mlifb, CCdflm, Uzd})
      6'd14: Mmiaej2 = 32'd2541311358 ^ 32'd2527372146;
      6'd39: Mmiaej2 = 32'd738229279 ^ 32'o34664350572 ^ 32'o35303055551;
      6'h1e: Mmiaej2 = 32'h63ca4b4 ^ 32'd1090138779 ^ 32'h471b6023;
      6'o62: Mmiaej2 = 32'd436547407 ^ 32'h19dffc7b ^ 32'b00000010000001110010010100111000;
      6'd2: Mmiaej2 = 32'b00000010100100111111001110011010 ^ 32'h34e0596;
      6'o35: Mmiaej2 = 32'o15101362425 ^ 32'o15066011431;
      6'd26: Mmiaej2 = 32'b11110001110001111000000000010000 ^ 32'h40f98c29 ^ 32'hb0e3fa35;
      6'h30: Mmiaej2 = 32'h5fd5fbb0 ^ 32'o13602006674;
      6'b001100: Mmiaej2 = 32'd176636439 ^ 32'o1326532033;
      6'd43: Mmiaej2 = 32'b10111111100001010110010010011010 ^ 32'o27626111226;
      6'o56: Mmiaej2 = 32'o24276103635 ^ 32'd2737140113;
      6'o75: Mmiaej2 = 32'b01011000110101010011110010001100 ^ 32'b01011001000010001100101010000000;
      6'o44: Mmiaej2 = 32'b11010000001011001000100000001010 ^ 32'd693376507 ^ 32'hf8a56bfd;
      6'd25: Mmiaej2 = 32'd1506198817 ^ 32'd462622806 ^ 32'h4388237b;
      6'd16: Mmiaej2 = 32'b10110010010101011001100000110110 ^ 32'hb3886e3a;
      6'b000101: Mmiaej2 = 32'b11101111100010100100001100000000 ^ 32'o30404715425 ^ 32'd709111321;
      6'b000011: Mmiaej2 = 32'o25450075454 ^ 32'o33337721656 ^ 32'd1979854478;
      6'h1b: Mmiaej2 = 32'b11111100000000111101100101000000 ^ 32'b00000001011001000001000010111011 ^ 32'b11111100101110100011111111110111;
      6'b110110: Mmiaej2 = 32'hc27cf35d ^ 32'd3282109777;
      6'b101010: Mmiaej2 = 32'o6141462030 ^ 32'b00110000010110111001001000010100;
      6'o76: Mmiaej2 = 32'h6e4b71f9 ^ 32'h6f9687f5;
      6'h11: Mmiaej2 = 32'o17141257050 ^ 32'h4b9a9bb7 ^ 32'd868365203;
      6'd24: Mmiaej2 = 32'hc11b0d40 ^ 32'o30061575514;
      6'o70: Mmiaej2 = 32'hb752dd98 ^ 32'd3062836116;
      6'h3a: Mmiaej2 = 32'b01100101101001111010011001100001 ^ 32'b01100100011110100101000001101101;
      6'h2c: Mmiaej2 = 32'b00011111011010110010001001100111 ^ 32'h1eb6d46b;
      6'b010011: Mmiaej2 = 32'h40a0faa4 ^ 32'h417d0ca8;
      6'o13: Mmiaej2 = 32'o1113420031 ^ 32'o1074753025;
      6'o42: Mmiaej2 = 32'o37451001200 ^ 32'o37536372214;
      6'b011111: Mmiaej2 = 32'h46f1a3ad ^ 32'o2340570650 ^ 32'd1420731401;
      6'b111111: Mmiaej2 = 32'o7335055634 ^ 32'b00111010101010011010110110010000;
      6'o34: Mmiaej2 = 32'o31133425453 ^ 32'hc8b3dd27;
      6'o71: Mmiaej2 = 32'o33015767545 ^ 32'b11011001111010100001100101101001;
      6'h0: Mmiaej2 = 32'h85ad1eec ^ 32'd3194900012 ^ 32'd975087308;
      6'h4: Mmiaej2 = 32'h8e1e0fae ^ 32'o20631711667 ^ 32'h9a46a15;
      6'hf: Mmiaej2 = 32'b00110010011001001110110011010111 ^ 32'b00110011101110010001101011011011;
      6'hd: Mmiaej2 = 32'b10000000010000010001101100000110 ^ 32'h93c2496a ^ 32'b00010010010111101010010001100000;
      6'h3c: Mmiaej2 = 32'hc4f0d7c9 ^ 32'o5564330713 ^ 32'he8fc900e;
      6'o1: Mmiaej2 = 32'd2544105416 ^ 32'd2524840388;
      6'o57: Mmiaej2 = 32'b10100110010000011010100101101101 ^ 32'b01110100111100100100111011111010 ^ 32'o32333410633;
      6'h23: Mmiaej2 = 32'o14025073066 ^ 32'b01100001100010011000000000111010;
      6'd33: Mmiaej2 = 32'hb99747b ^ 32'o1221101167;
      6'h34: Mmiaej2 = 32'o10502765620 ^ 32'h44d61d9c;
      6'd18: Mmiaej2 = 32'b11001111010010001001000001011010 ^ 32'b11001110100101010110011001010110;
      6'b110101: Mmiaej2 = 32'o11055064577 ^ 32'o11132317563;
      6'd41: Mmiaej2 = 32'b10101110010000011101100001111100 ^ 32'hceb9fb97 ^ 32'b01100001001001011101010111100111;
      6'd45: Mmiaej2 = 32'b11000110100101011111010011000100 ^ 32'o12640715640 ^ 32'h91cb9968;
      6'o12: Mmiaej2 = 32'h71d5ce1c ^ 32'd557584257 ^ 32'd1362376593;
      6'o61: Mmiaej2 = 32'o35727172462 ^ 32'o640030513 ^ 32'd3892392565;
      6'b111011: Mmiaej2 = 32'b01000111101001100101000001100000 ^ 32'b01000001000011011101111100110110 ^ 32'o735474532;
      6'b100101: Mmiaej2 = 32'o21476112170 ^ 32'o25345100601 ^ 32'd649192437;
      6'h26: Mmiaej2 = 32'b01110111101111110011110110001001 ^ 32'd1986186117;
      6'b100000: Mmiaej2 = 32'b10101011101011001101000111011100 ^ 32'd2690664351 ^ 32'o1204260117;
      6'd20: Mmiaej2 = 32'o37552471256 ^ 32'hce1ccdf9 ^ 32'b00110010011010110100100101011011;
      6'h8: Mmiaej2 = 32'o15116130215 ^ 32'h68e54681;
      6'b001001: Mmiaej2 = 32'h16ae88fb ^ 32'hdaa95bef ^ 32'd3453625624;
      6'b101000: Mmiaej2 = 32'b00001110110010101100000101010110 ^ 32'b00001111000101110011011101011010;
      6'o6: Mmiaej2 = 32'o31706370756 ^ 32'b11001110110001000000011111100010;
      6'b110011: Mmiaej2 = 32'o1325276447 ^ 32'b00001010100010001000101100101011;
      6'd7: Mmiaej2 = 32'o26543236710 ^ 32'h9450cbc4;
      6'd23: Mmiaej2 = 32'b11110000000011011100000110011110 ^ 32'b11011000000100011100010110011010 ^ 32'b00001001110000011111001000001000;
      6'h16: Mmiaej2 = 32'd264944835 ^ 32'd236407503;
      6'h37: Mmiaej2 = 32'h946bf491 ^ 32'b01100001000101110110100000010010 ^ 32'd3567348367;
      6'd21: Mmiaej2 = 32'h317d6249 ^ 32'b00110000101000001001010001000101;

      default: Mmiaej2 = 32'hdead_dead;
    endcase
  end

  logic [7:0] pFiH5vTGl;
  assign pFiH5vTGl = ra2VgcBEzc[7:0];

  always_ff @(posedge clk_i) begin
    if(rst_i) begin
      data <= '0;
    end
    else if (gUruyn1hzjChHha47v[32'o5102152502 ^ 32'o5102152500]) begin
      data <= '0;
    end
    else if(Mmiaej2[32'h5173ee4c ^ 32'o12134767121]) begin
      data <= pFiH5vTGl;
    end
    else begin
      data <= data;
    end
  end
  assign CCdflm = Y2pd == (32'h4300c627 ^ 32'h1eac865e ^ 32'b01011101101011000100000001111001);

  logic tzBmaC;
  logic [31:0] Ms1Hk7Iek2EKZQuQME347y;
  always_comb begin
    case ({YAhtnxC5bxEVGCn, Uzd, cWdgq, parity_en, B4zEGLaAwyO6, Gdxya89mlifb})
      6'b001101: Ms1Hk7Iek2EKZQuQME347y = 32'o33751265117 ^ 32'd3613260120;
      6'o13: Ms1Hk7Iek2EKZQuQME347y = 32'd4137752744 ^ 32'o37163167253 ^ 32'd127231252;
      6'b110010: Ms1Hk7Iek2EKZQuQME347y = 32'd4189286840 ^ 32'd2439194499 ^ 32'h6028c52c;
      6'd9: Ms1Hk7Iek2EKZQuQME347y = 32'o35353211177 ^ 32'o17120402427 ^ 32'o23205702177;
      6'd63: Ms1Hk7Iek2EKZQuQME347y = 32'b00101111111010010100100011110111 ^ 32'h2713dbe0;
      6'o4: Ms1Hk7Iek2EKZQuQME347y = 32'o13360237053 ^ 32'h5339ad3c;
      6'b000001: Ms1Hk7Iek2EKZQuQME347y = 32'o32251270643 ^ 32'o33227361264;
      6'o35: Ms1Hk7Iek2EKZQuQME347y = 32'hc88eece7 ^ 32'd3228991472;
      6'b010101: Ms1Hk7Iek2EKZQuQME347y = 32'o36152502530 ^ 32'd4182906447;
      6'b101010: Ms1Hk7Iek2EKZQuQME347y = 32'b11111101010010011110110100100110 ^ 32'b00100000010011100000111001100000 ^ 32'b11010101111111110111000001010001;
      6'b101011: Ms1Hk7Iek2EKZQuQME347y = 32'd3715952943 ^ 32'hd5846238;
      6'o7: Ms1Hk7Iek2EKZQuQME347y = 32'd1215726386 ^ 32'h52993c0 ^ 32'd1168606181;
      6'h12: Ms1Hk7Iek2EKZQuQME347y = 32'd1109369178 ^ 32'd1470538531 ^ 32'o3520310556;
      6'o37: Ms1Hk7Iek2EKZQuQME347y = 32'h63d55ec5 ^ 32'h5652ef65 ^ 32'd1031742135;
      6'h28: Ms1Hk7Iek2EKZQuQME347y = 32'h818375c3 ^ 32'o13531511200 ^ 32'o32407272124;
      6'o6: Ms1Hk7Iek2EKZQuQME347y = 32'o127264611 ^ 32'o34557557441 ^ 32'b11101100000110110010010110111111;
      6'hf: Ms1Hk7Iek2EKZQuQME347y = 32'd61230081 ^ 32'o1327557426;
      6'b100001: Ms1Hk7Iek2EKZQuQME347y = 32'b00001110110111011101100110000001 ^ 32'h6254a96;
      6'b110101: Ms1Hk7Iek2EKZQuQME347y = 32'o22667266123 ^ 32'd2653290308;
      6'd36: Ms1Hk7Iek2EKZQuQME347y = 32'b10101001011101101111101111011111 ^ 32'ha18e68c8;
      6'd45: Ms1Hk7Iek2EKZQuQME347y = 32'b01110100010110011110111000001101 ^ 32'd2090958106;
      6'b100010: Ms1Hk7Iek2EKZQuQME347y = 32'b10010011111101010111001111000110 ^ 32'd79399243 ^ 32'h9fb6699a;
      6'o10: Ms1Hk7Iek2EKZQuQME347y = 32'b10101111100010100101001100011111 ^ 32'b10100111011100101100000000001000;
      6'o70: Ms1Hk7Iek2EKZQuQME347y = 32'h4b7e1eb2 ^ 32'hcf31a079 ^ 32'b10001100101101110010110111011100;
      6'd54: Ms1Hk7Iek2EKZQuQME347y = 32'h3eae9733 ^ 32'o14127351641 ^ 32'b01010111000010111101011110000101;
      6'b000011: Ms1Hk7Iek2EKZQuQME347y = 32'b00101011001100011101110010110011 ^ 32'b01101100111111110001110111000000 ^ 32'b01001111001101100101001001100100;
      6'd35: Ms1Hk7Iek2EKZQuQME347y = 32'd1097232383 ^ 32'hc062c0f1 ^ 32'h89fc3c19;
      6'o57: Ms1Hk7Iek2EKZQuQME347y = 32'h8549c521 ^ 32'd2377209398;
      6'o61: Ms1Hk7Iek2EKZQuQME347y = 32'd3369499619 ^ 32'hefbb5416 ^ 32'h2f95bce2;
      6'b010100: Ms1Hk7Iek2EKZQuQME347y = 32'b00110001010110000000101000011010 ^ 32'h39a0990d;
      6'h13: Ms1Hk7Iek2EKZQuQME347y = 32'o5433110322 ^ 32'o23463122620 ^ 32'o27026123125;
      6'o16: Ms1Hk7Iek2EKZQuQME347y = 32'o5723225300 ^ 32'o4755334727;
      6'b001010: Ms1Hk7Iek2EKZQuQME347y = 32'h68d09613 ^ 32'd525324673 ^ 32'h7f67d485;
      6'o47: Ms1Hk7Iek2EKZQuQME347y = 32'o37610656050 ^ 32'b11110110110110111100111100111111;
      6'o2: Ms1Hk7Iek2EKZQuQME347y = 32'he5c49f5d ^ 32'b10111110010000011001001011011110 ^ 32'o12337317224;
      6'd57: Ms1Hk7Iek2EKZQuQME347y = 32'o23143462273 ^ 32'd2440492972;
      6'h34: Ms1Hk7Iek2EKZQuQME347y = 32'd2761539638 ^ 32'd2486762226 ^ 32'b00111000010110011010100111010011;
      6'o30: Ms1Hk7Iek2EKZQuQME347y = 32'o14306066724 ^ 32'b00011011001011001000011011010110 ^ 32'b01110000110011000111100000010101;
      6'h19: Ms1Hk7Iek2EKZQuQME347y = 32'o4060712276 ^ 32'd393487292 ^ 32'd1062151189;
      6'h1a: Ms1Hk7Iek2EKZQuQME347y = 32'd1662721241 ^ 32'd1810075598;
      6'o21: Ms1Hk7Iek2EKZQuQME347y = 32'hba0c63c6 ^ 32'b10110010111101001111000011010001;
      6'o45: Ms1Hk7Iek2EKZQuQME347y = 32'o15354465702 ^ 32'd4194278056 ^ 32'h9ab5627d;
      6'h33: Ms1Hk7Iek2EKZQuQME347y = 32'b01011011100101100110101111010001 ^ 32'd3392120704 ^ 32'b10011001010000110101111101000110;
      6'o56: Ms1Hk7Iek2EKZQuQME347y = 32'b01111010001101001111110110011100 ^ 32'h72cc6e8b;
      6'b111110: Ms1Hk7Iek2EKZQuQME347y = 32'd1572344914 ^ 32'd4080805520 ^ 32'd2793185749;
      6'b001100: Ms1Hk7Iek2EKZQuQME347y = 32'b11100010000011010100101000100011 ^ 32'd3941980468;
      6'o72: Ms1Hk7Iek2EKZQuQME347y = 32'h16262545 ^ 32'o3667533122;
      6'o36: Ms1Hk7Iek2EKZQuQME347y = 32'o30642111122 ^ 32'o37775175540 ^ 32'b00110001100001001111101000100101;
      6'h0: Ms1Hk7Iek2EKZQuQME347y = 32'd3969910535 ^ 32'o34426112020;
      6'd22: Ms1Hk7Iek2EKZQuQME347y = 32'o7343571445 ^ 32'o6335460062;
      6'h1c: Ms1Hk7Iek2EKZQuQME347y = 32'o27374776115 ^ 32'hb30b6f5a;
      6'o74: Ms1Hk7Iek2EKZQuQME347y = 32'b00100011010001101101011100010000 ^ 32'b00101011101111100100010000000111;
      6'o33: Ms1Hk7Iek2EKZQuQME347y = 32'o7337760421 ^ 32'heffa8aad ^ 32'b11011100011111011111100010101011;
      6'b111011: Ms1Hk7Iek2EKZQuQME347y = 32'o23037130714 ^ 32'd3932785086 ^ 32'b01111010111011111010101101100101;
      6'o46: Ms1Hk7Iek2EKZQuQME347y = 32'd3186732344 ^ 32'hdde151a0 ^ 32'b01101000111010000110111110001111;
      6'o67: Ms1Hk7Iek2EKZQuQME347y = 32'o33403710247 ^ 32'hd4f503b0;
      6'h29: Ms1Hk7Iek2EKZQuQME347y = 32'b00110011000110001001110011001100 ^ 32'b00111011111000000000111111011011;
      6'd5: Ms1Hk7Iek2EKZQuQME347y = 32'd1358988791 ^ 32'd3300201142 ^ 32'o23523202126;
      6'd44: Ms1Hk7Iek2EKZQuQME347y = 32'b11011111010110110110101100001100 ^ 32'd3743037766 ^ 32'd146391389;
      6'o40: Ms1Hk7Iek2EKZQuQME347y = 32'd2436372111 ^ 32'o22257126063 ^ 32'hb7c29ab;
      6'o20: Ms1Hk7Iek2EKZQuQME347y = 32'b01111011001101001100111110111111 ^ 32'o11350172673 ^ 32'o7033124423;
      6'h17: Ms1Hk7Iek2EKZQuQME347y = 32'o17703170211 ^ 32'o16775061636;
      6'h30: Ms1Hk7Iek2EKZQuQME347y = 32'heac0384f ^ 32'o26105346401 ^ 32'h532d6659;
      6'b111101: Ms1Hk7Iek2EKZQuQME347y = 32'h8e0a8415 ^ 32'd2264012546;
      default: Ms1Hk7Iek2EKZQuQME347y = 32'hdead_dead;
    endcase
  end

  logic [31:0] N70LunC3adr;
  always_comb begin
    case ({YAhtnxC5bxEVGCn, parity_en, busy, Gdxya89mlifb, Uzd, tzBmaC})
      6'd51: N70LunC3adr = 32'o2617214770 ^ 32'b01100011111101111000101100110001;
      6'd30: N70LunC3adr = 32'hcc273787 ^ 32'b10111001111011011010010101001110;
      6'o41: N70LunC3adr = 32'd3442781752 ^ 32'o27077436361;
      6'h19: N70LunC3adr = 32'o21657165761 ^ 32'd3639197280 ^ 32'o4347743530;
      6'o72: N70LunC3adr = 32'h56a9b6c5 ^ 32'b00100011011000110010010000001100;
      6'h2f: N70LunC3adr = 32'b00000010001000101011001101011101 ^ 32'b01110111111010010010000110010100;
      6'h9: N70LunC3adr = 32'd3919098990 ^ 32'o23424423247;
      6'b010011: N70LunC3adr = 32'o25706037655 ^ 32'b11101110110101111110100101101110 ^ 32'o6401242012;
      6'b110000: N70LunC3adr = 32'had3371d8 ^ 32'd1171831056 ^ 32'd2636208641;
      6'b010000: N70LunC3adr = 32'd3630077391 ^ 32'd4106048578 ^ 32'd1495880516;
      6'b001101: N70LunC3adr = 32'ha93945e5 ^ 32'd3706967852;
      6'h32: N70LunC3adr = 32'b01101011000100000001100010001000 ^ 32'hafc13153 ^ 32'd2971384594;
      6'b010111: N70LunC3adr = 32'b10100010000001110110001000101101 ^ 32'd647163765 ^ 32'o36127417621;
      6'he: N70LunC3adr = 32'hb77f43f0 ^ 32'd3266695481;
      6'o35: N70LunC3adr = 32'o30521075135 ^ 32'b10110000100011101110100010010100;
      6'h3e: N70LunC3adr = 32'hb0fa72ac ^ 32'hc530e065;
      6'h20: N70LunC3adr = 32'h8d544b19 ^ 32'd2331862750 ^ 32'b01110010011000111011111100001110;
      6'o6: N70LunC3adr = 32'b10101100010101010101101110001100 ^ 32'b11011001100111111100100101000101;
      6'h0: N70LunC3adr = 32'o27544637554 ^ 32'd449366871 ^ 32'b11010010100100010110011011110010;
      6'o1: N70LunC3adr = 32'd1391804490 ^ 32'o24614313474 ^ 32'h810e45bf;
      6'b110110: N70LunC3adr = 32'd3431120193 ^ 32'h82fdd87 ^ 32'hb167f20f;
      6'd39: N70LunC3adr = 32'hc7f676ca ^ 32'hec5d5861 ^ 32'o13630136142;
      6'd12: N70LunC3adr = 32'd3198228442 ^ 32'hcb6b8513;
      6'h8: N70LunC3adr = 32'b01111111100100001111110000000010 ^ 32'ha5a6ecb;
      6'b100011: N70LunC3adr = 32'h9f6d0c7a ^ 32'o24602736240 ^ 32'b01001100101011000010001000010011;
      6'b110111: N70LunC3adr = 32'he7d0d521 ^ 32'hbebb92b3 ^ 32'o5450152533;
      6'o55: N70LunC3adr = 32'b01000101111111001001010101011000 ^ 32'o15121511031 ^ 32'b01011001011100001001010110001000;
      6'b101011: N70LunC3adr = 32'hd5099c82 ^ 32'b10100000110000110000111001001011;
      6'b000011: N70LunC3adr = 32'd2797617917 ^ 32'b11110101101110000000101010000000 ^ 32'b00100110101100101101101010110100;
      6'd28: N70LunC3adr = 32'hf41ddb43 ^ 32'o20165644612;
      6'd17: N70LunC3adr = 32'b01001010010011110010101001110000 ^ 32'o7741334271;
      6'd22: N70LunC3adr = 32'h63261ec7 ^ 32'd384601102;
      6'h3c: N70LunC3adr = 32'hbffd22e8 ^ 32'd3392647201;
      6'o70: N70LunC3adr = 32'o24273550365 ^ 32'd3609477692;
      6'b010100: N70LunC3adr = 32'ha50064c7 ^ 32'd3502962190;
      6'h26: N70LunC3adr = 32'd1634415701 ^ 32'd346138268;
      6'h2e: N70LunC3adr = 32'o7165325552 ^ 32'h4c1f39a3;
      6'b111101: N70LunC3adr = 32'hf33f33ce ^ 32'd2601140310 ^ 32'h1dffe151;
      6'h3b: N70LunC3adr = 32'h298aed3d ^ 32'h2dd8046d ^ 32'd1905818521;
      6'b011010: N70LunC3adr = 32'o16121007371 ^ 32'o3376022737 ^ 32'd527874543;
      6'o5: N70LunC3adr = 32'b10100001101111100010011000000000 ^ 32'o10517031350 ^ 32'b10010001010010001000011000100001;
      6'h2a: N70LunC3adr = 32'ha1b63a4b ^ 32'b01111100000011100101010110100100 ^ 32'o25034576446;
      6'h4: N70LunC3adr = 32'b10001010101011100011001110101001 ^ 32'o32626044416 ^ 32'o5117164156;
      6'h3f: N70LunC3adr = 32'h695ad93 ^ 32'b01110011010111100011111101011010;
      6'd24: N70LunC3adr = 32'd3227822064 ^ 32'd2878952916 ^ 32'h1e3760ed;
      6'b011011: N70LunC3adr = 32'b10110000101011001110101111100110 ^ 32'o6120640113 ^ 32'hf4253964;
      6'o25: N70LunC3adr = 32'hc9f0946d ^ 32'b10000001110010100100110001001100 ^ 32'b00111101111100000100101011101000;
      6'd31: N70LunC3adr = 32'd4102483061 ^ 32'd1494636789 ^ 32'd3629852233;
      6'b110001: N70LunC3adr = 32'd2469654835 ^ 32'o34676261772;
      6'h34: N70LunC3adr = 32'd2149109622 ^ 32'b11110101110100100101110110111111;
      6'o13: N70LunC3adr = 32'hcc53352e ^ 32'h14258722 ^ 32'hadbc20c5;
      6'b001111: N70LunC3adr = 32'o21117752577 ^ 32'h17c5a3ab ^ 32'o35314362035;
      6'h29: N70LunC3adr = 32'h3a7aa2c2 ^ 32'h4fb0300b;
      6'b111001: N70LunC3adr = 32'o2062162745 ^ 32'ha651f7ee ^ 32'o30324700302;
      6'ha: N70LunC3adr = 32'b11101000101100101101111110000110 ^ 32'b10011101011110000100110101001111;
      6'b100101: N70LunC3adr = 32'hb5a1c9bb ^ 32'd2598522145 ^ 32'o13242213123;
      6'h2: N70LunC3adr = 32'd602465650 ^ 32'h848331d6 ^ 32'hd2a1466d;
      6'h35: N70LunC3adr = 32'o16325017771 ^ 32'd111054128;
      6'd7: N70LunC3adr = 32'b01000000011000011101001000101001 ^ 32'd900350176;
      6'b100010: N70LunC3adr = 32'hb28fc09c ^ 32'hc7455255;
      6'd40: N70LunC3adr = 32'heed249fb ^ 32'o23306155462;
      6'd44: N70LunC3adr = 32'he9140290 ^ 32'o23467510131;
      6'd18: N70LunC3adr = 32'd3548819580 ^ 32'd2790007477;
      6'h24: N70LunC3adr = 32'hf066528d ^ 32'd2242691140;
      default: N70LunC3adr = 32'hdead_dead;
    endcase
  end

  logic [16:0] sdCSHTFRGa6pA;
  assign sdCSHTFRGa6pA = ra2VgcBEzc[16:0];

  always_ff @(posedge clk_i) begin
    if(rst_i) begin
      baudrate <= 9600;
    end
    else if (Ms1Hk7Iek2EKZQuQME347y[32'o34423457114 ^ 32'o34423457135]) begin
      baudrate <= 9600;
    end
    else if(N70LunC3adr[32'h2aa8fa8 ^ 32'h280bf186 ^ 32'b00101010101000010111111000111110]) begin
      baudrate <= sdCSHTFRGa6pA;
    end
    else begin
      baudrate <= baudrate;
    end
  end

  logic lYDnXNr;
  assign lYDnXNr = (Y2pd == (32'o5304103005 ^ 32'o21020144777 ^ 32'ha3504fea));
  logic [31:0] EbCa5mgVyDjWmA;

  always_comb begin
    case ({YAhtnxC5bxEVGCn, lYDnXNr, parity_en, Uzd, B4zEGLaAwyO6, Gdxya89mlifb, ra2VgcBEzc[0]})
      7'o22: EbCa5mgVyDjWmA = 32'o132064763 ^ 32'h3f79ae32 ^ 32'h55806141;
      7'b0100011: EbCa5mgVyDjWmA = 32'o3574452700 ^ 32'b01110110011000111111011101000000;
      7'd23: EbCa5mgVyDjWmA = 32'd1057395459 ^ 32'h54973583;
      7'o76: EbCa5mgVyDjWmA = 32'o27023672617 ^ 32'd1391854611 ^ 32'h8128d31c;
      7'o7: EbCa5mgVyDjWmA = 32'b11010101010101110001101001011001 ^ 32'hbec6b8d9;
      7'b1010001: EbCa5mgVyDjWmA = 32'd1871413174 ^ 32'o34565033541 ^ 32'b11100001110011101110111001010111;
      7'o74: EbCa5mgVyDjWmA = 32'h68bef637 ^ 32'd3642659718 ^ 32'o33214341461;
      7'o151: EbCa5mgVyDjWmA = 32'o404765352 ^ 32'd1870809194;
      7'b1100011: EbCa5mgVyDjWmA = 32'h59c0867 ^ 32'd1735843965 ^ 32'o1136645232;
      7'o122: EbCa5mgVyDjWmA = 32'o16011650615 ^ 32'd464975629;
      7'd126: EbCa5mgVyDjWmA = 32'd3875967112 ^ 32'o21445631010;
      7'o63: EbCa5mgVyDjWmA = 32'd3001622358 ^ 32'o33136134726;
      7'd76: EbCa5mgVyDjWmA = 32'h92f832b7 ^ 32'b11111001011010011001000000110111;
      7'd90: EbCa5mgVyDjWmA = 32'had986f4e ^ 32'd3322530254;
      7'd0: EbCa5mgVyDjWmA = 32'd3812247673 ^ 32'd2292968185;
      7'ha: EbCa5mgVyDjWmA = 32'b10010010101110000011110001110010 ^ 32'd4180254450;
      7'd17: EbCa5mgVyDjWmA = 32'b10100001000011010100111110101101 ^ 32'o35051610563 ^ 32'b00100010001110111111100001011110;
      7'h6a: EbCa5mgVyDjWmA = 32'h8e209a0 ^ 32'hb1fd252a ^ 32'b11010010100011101000111000001010;
      7'd29: EbCa5mgVyDjWmA = 32'o11740617531 ^ 32'o4404534731;
      7'b0110110: EbCa5mgVyDjWmA = 32'o7627522332 ^ 32'd16044852 ^ 32'b01010101001110111101000101101110;
      7'h49: EbCa5mgVyDjWmA = 32'o36206126651 ^ 32'h99890f29;
      7'd61: EbCa5mgVyDjWmA = 32'hf0662844 ^ 32'o14766771467 ^ 32'hfc2c7df3;
      7'b1111100: EbCa5mgVyDjWmA = 32'o3521530165 ^ 32'b01110110110101110001011011110101;
      7'b1010011: EbCa5mgVyDjWmA = 32'b00001110010101111011110011011111 ^ 32'o14561415137;
      7'o163: EbCa5mgVyDjWmA = 32'b00010001111111000100010110010001 ^ 32'h7a6de311;
      7'd21: EbCa5mgVyDjWmA = 32'b00101010101010100101000111111000 ^ 32'b10101000110011001000001101101010 ^ 32'he9f77412;
      7'o20: EbCa5mgVyDjWmA = 32'o37600775774 ^ 32'b11011100010000110001010001111010 ^ 32'd1238452486;
      7'd34: EbCa5mgVyDjWmA = 32'o37754747625 ^ 32'he8b4c5d6 ^ 32'd2090248387;
      7'b1000110: EbCa5mgVyDjWmA = 32'o1427627533 ^ 32'd1884362349 ^ 32'o2747715666;
      7'd98: EbCa5mgVyDjWmA = 32'b01010101000010001000101100001001 ^ 32'o7646224611;
      7'b0111000: EbCa5mgVyDjWmA = 32'h64557702 ^ 32'd3467552707 ^ 32'b11000001011010100111011001000001;
      7'h78: EbCa5mgVyDjWmA = 32'hef35525a ^ 32'b10000100101001001111010011011010;
      7'o116: EbCa5mgVyDjWmA = 32'd3742197671 ^ 32'o20771671135 ^ 32'o6336733572;
      7'o45: EbCa5mgVyDjWmA = 32'hab1563ee ^ 32'hc084c16e;
      7'hf: EbCa5mgVyDjWmA = 32'd1017579748 ^ 32'b01010111001101101010101001100100;
      7'd32: EbCa5mgVyDjWmA = 32'o14407022107 ^ 32'hf8d86c7;
      7'o57: EbCa5mgVyDjWmA = 32'h27530fe8 ^ 32'd1287825768;
      7'o140: EbCa5mgVyDjWmA = 32'b10001101100011110101110110011001 ^ 32'o21175442155 ^ 32'o15772135564;
      7'h5f: EbCa5mgVyDjWmA = 32'h5cac8f0d ^ 32'o6717226615;
      7'd64: EbCa5mgVyDjWmA = 32'h2b319f8c ^ 32'hbeebb58e ^ 32'b11111110010010111000100010000010;
      7'd48: EbCa5mgVyDjWmA = 32'o2570322332 ^ 32'b10010111111111100111111110001000 ^ 32'b11101001100011100111110111010010;
      7'b1110100: EbCa5mgVyDjWmA = 32'o31002304640 ^ 32'b10100011100110000010111100100000;
      7'b1000111: EbCa5mgVyDjWmA = 32'o26446210446 ^ 32'h99f17411 ^ 32'd1190774711;
      7'b1101100: EbCa5mgVyDjWmA = 32'b00001100101001000101000100000010 ^ 32'd2669964437 ^ 32'hf8119f17;
      7'o73: EbCa5mgVyDjWmA = 32'b00101100111000011110000111101100 ^ 32'h4770476c;
      7'o33: EbCa5mgVyDjWmA = 32'd1598780250 ^ 32'd139131655 ^ 32'b00111100100100000010111011011101;
      7'b0001000: EbCa5mgVyDjWmA = 32'o761575714 ^ 32'o15425654514;
      7'b1110010: EbCa5mgVyDjWmA = 32'h74e5538a ^ 32'o3735172412;
      7'o104: EbCa5mgVyDjWmA = 32'o444614032 ^ 32'o27652741272 ^ 32'd3517544480;
      7'd74: EbCa5mgVyDjWmA = 32'd3547333056 ^ 32'ha56a8c1f ^ 32'd495660895;
      7'h65: EbCa5mgVyDjWmA = 32'b00101011000001101011000101111001 ^ 32'h409713f9;
      7'h13: EbCa5mgVyDjWmA = 32'd723664635 ^ 32'o35146162527 ^ 32'd2838199596;
      7'd89: EbCa5mgVyDjWmA = 32'o32610505275 ^ 32'h4d30f7a5 ^ 32'o36040755630;
      7'h7d: EbCa5mgVyDjWmA = 32'he9972542 ^ 32'ha954b6b8 ^ 32'b00101011010100100011010101111010;
      7'd50: EbCa5mgVyDjWmA = 32'o22531053165 ^ 32'hfef5f0f5;
      7'b1101011: EbCa5mgVyDjWmA = 32'h91503ca6 ^ 32'b11101111010101001001010100000100 ^ 32'b00010101100101010000111100100010;
      7'h55: EbCa5mgVyDjWmA = 32'b00011111100001111011011110001111 ^ 32'd1947603215;
      7'he: EbCa5mgVyDjWmA = 32'd3562969044 ^ 32'd2188800996 ^ 32'd1035552432;
      7'hd: EbCa5mgVyDjWmA = 32'b01110100001010100110010100100110 ^ 32'd3308037185 ^ 32'o33245661747;
      7'b1011101: EbCa5mgVyDjWmA = 32'he75fd828 ^ 32'o21463477250;
      7'h5: EbCa5mgVyDjWmA = 32'd2345549419 ^ 32'd3764362475;
      7'h45: EbCa5mgVyDjWmA = 32'd976999875 ^ 32'h51aa7743;
      7'h5c: EbCa5mgVyDjWmA = 32'd25584060 ^ 32'd3278773428 ^ 32'd2843335560;
      7'o171: EbCa5mgVyDjWmA = 32'd3778413982 ^ 32'd2326242078;
      7'd57: EbCa5mgVyDjWmA = 32'h389595c0 ^ 32'o37215521117 ^ 32'b10101001001100101001000100001111;
      7'd12: EbCa5mgVyDjWmA = 32'h8cd802c9 ^ 32'o6152237477 ^ 32'b11010110111000001001111101110110;
      7'h6d: EbCa5mgVyDjWmA = 32'hf8273d47 ^ 32'd5712625 ^ 32'b10010011111000011011010100110110;
      7'b1101111: EbCa5mgVyDjWmA = 32'd2255462157 ^ 32'b11110001010101011001111111110011 ^ 32'o3452721176;
      7'o3: EbCa5mgVyDjWmA = 32'o2513673212 ^ 32'hbd65e872 ^ 32'd3285924984;
      7'o30: EbCa5mgVyDjWmA = 32'b01100011111010010100010011110010 ^ 32'h878e272;
      7'd86: EbCa5mgVyDjWmA = 32'b01110010011000100110000101011000 ^ 32'd435406808;
      7'b0011001: EbCa5mgVyDjWmA = 32'd1069586730 ^ 32'o31156772761 ^ 32'd2649410139;
      7'b1100111: EbCa5mgVyDjWmA = 32'd2489104982 ^ 32'd751176986 ^ 32'o32302612714;
      7'b1010111: EbCa5mgVyDjWmA = 32'o126315027 ^ 32'h4e97f187 ^ 32'b00100100010111111100110100010000;
      7'h1f: EbCa5mgVyDjWmA = 32'b00000100001011011010110111110101 ^ 32'b01110111100000111111101000111100 ^ 32'd406843721;
      7'o36: EbCa5mgVyDjWmA = 32'b10100001000101000000000000011000 ^ 32'hca85a698;
      7'h37: EbCa5mgVyDjWmA = 32'd505568303 ^ 32'h75b3faaf;
      7'h50: EbCa5mgVyDjWmA = 32'b00011001100110100001000000110010 ^ 32'h720bb6b2;
      7'h2a: EbCa5mgVyDjWmA = 32'b10001111111111110101111110111001 ^ 32'o26744073457 ^ 32'o12377505026;
      7'o130: EbCa5mgVyDjWmA = 32'o2744234645 ^ 32'o7555112050 ^ 32'o10155005415;
      7'd67: EbCa5mgVyDjWmA = 32'o17510766615 ^ 32'o2654447415;
      7'o136: EbCa5mgVyDjWmA = 32'o6247070360 ^ 32'o11044513200 ^ 32'h119f44f0;
      7'b0101100: EbCa5mgVyDjWmA = 32'o10264236616 ^ 32'b00101001010000001001111100001110;
      7'o172: EbCa5mgVyDjWmA = 32'h7fc97415 ^ 32'o14702254430 ^ 32'd1934725005;
      7'h21: EbCa5mgVyDjWmA = 32'd588863211 ^ 32'b00001100001010111010101100110100 ^ 32'd1151557471;
      7'd97: EbCa5mgVyDjWmA = 32'd381929066 ^ 32'b01111101010100100110010011101010;
      7'o101: EbCa5mgVyDjWmA = 32'd2616857153 ^ 32'hf06bb0c1;
      7'b0110001: EbCa5mgVyDjWmA = 32'b10111101000100010110111111111000 ^ 32'd627651425 ^ 32'b11110011111010011111101000011001;
      7'h6e: EbCa5mgVyDjWmA = 32'd1712015651 ^ 32'hd9aeba3;
      7'o110: EbCa5mgVyDjWmA = 32'd4042923948 ^ 32'b10011011011010111011110100101100;
      7'b1110110: EbCa5mgVyDjWmA = 32'h8b6c6095 ^ 32'd3774727701;
      7'h4b: EbCa5mgVyDjWmA = 32'd1999785610 ^ 32'b00011100101000111110110000001010;
      7'h9: EbCa5mgVyDjWmA = 32'h19913ce8 ^ 32'o26217602530 ^ 32'hc03f9b30;
      7'o55: EbCa5mgVyDjWmA = 32'o25572326407 ^ 32'd4203183826 ^ 32'h3cff7155;
      7'b1111011: EbCa5mgVyDjWmA = 32'hcdeb7b36 ^ 32'b10100110011110101101110110110110;
      7'o44: EbCa5mgVyDjWmA = 32'b00011100011100011000111000111000 ^ 32'o31327675522 ^ 32'd3166656490;
      7'b0011100: EbCa5mgVyDjWmA = 32'o27611156240 ^ 32'b11110000001110111110011001010010 ^ 32'b00100101100011101001110001110010;
      7'b0000100: EbCa5mgVyDjWmA = 32'h8ee0f871 ^ 32'o34470436432 ^ 32'd26437611;
      7'd20: EbCa5mgVyDjWmA = 32'o25314126562 ^ 32'o30050205762;
      7'd63: EbCa5mgVyDjWmA = 32'd2120804695 ^ 32'h15f94fd7;
      7'h54: EbCa5mgVyDjWmA = 32'd2406027726 ^ 32'b11100100111110001011011101001110;
      7'd43: EbCa5mgVyDjWmA = 32'o12332513743 ^ 32'h15832eb1 ^ 32'd762847186;
      7'b0110101: EbCa5mgVyDjWmA = 32'd3841721351 ^ 32'o21010014364 ^ 32'b00000111010011011011101001110011;
      7'd39: EbCa5mgVyDjWmA = 32'b11100101000110010011100001100010 ^ 32'h8e889ae2;
      7'b0001011: EbCa5mgVyDjWmA = 32'h909c2c ^ 32'd1429848286 ^ 32'o7616177162;
      7'h4d: EbCa5mgVyDjWmA = 32'b11100100111101010000000111000111 ^ 32'o34326005561 ^ 32'o15417124066;
      7'o56: EbCa5mgVyDjWmA = 32'o10523640623 ^ 32'h2edee313;
      7'b1001111: EbCa5mgVyDjWmA = 32'd2199698873 ^ 32'd1880109399 ^ 32'b10011000100111010010111001101110;
      7'd52: EbCa5mgVyDjWmA = 32'h91ce02d4 ^ 32'b10011111101010110110001111110010 ^ 32'o14575143646;
      7'd102: EbCa5mgVyDjWmA = 32'd3030320578 ^ 32'hdf0ea742;
      7'd119: EbCa5mgVyDjWmA = 32'o10061052434 ^ 32'hb968c9f1 ^ 32'h923d3a6d;
      7'h5b: EbCa5mgVyDjWmA = 32'h3c3e461 ^ 32'd1750221537;
      7'd127: EbCa5mgVyDjWmA = 32'd4213818314 ^ 32'b11110000011101101000001001011111 ^ 32'b01100000110011101110001100010101;
      7'o161: EbCa5mgVyDjWmA = 32'b11100011001011110101001010010001 ^ 32'h2704c7ec ^ 32'b10101111101110100011001111111101;
      7'b0000001: EbCa5mgVyDjWmA = 32'h300df43b ^ 32'o33225337752 ^ 32'h81c9e951;
      7'b0011010: EbCa5mgVyDjWmA = 32'd985387451 ^ 32'o12112473473;
      7'd41: EbCa5mgVyDjWmA = 32'o32044377757 ^ 32'd502406741 ^ 32'b10100110111100100100001100111010;
      7'o72: EbCa5mgVyDjWmA = 32'h6d98a8ca ^ 32'd101255754;
      7'd38: EbCa5mgVyDjWmA = 32'b10000110110000100100101011111010 ^ 32'o35524764172;
      7'h70: EbCa5mgVyDjWmA = 32'd3245086081 ^ 32'b10101010111111011011001100000001;
      7'h6: EbCa5mgVyDjWmA = 32'd2924711768 ^ 32'b11000101110000100010110111011000;
      7'b1100100: EbCa5mgVyDjWmA = 32'd1060479763 ^ 32'o12451000623;
      7'b0010110: EbCa5mgVyDjWmA = 32'o17526102700 ^ 32'b10101110111110011101110100110010 ^ 32'b10111000001100001111111001110010;
      7'o102: EbCa5mgVyDjWmA = 32'o16461006026 ^ 32'b11110011001110010001110011110001 ^ 32'o35433131147;
      7'o50: EbCa5mgVyDjWmA = 32'b10011110010010100010101010000110 ^ 32'o36566704006;
      7'b1110101: EbCa5mgVyDjWmA = 32'ha34897e2 ^ 32'hc8d93162;
      7'o2: EbCa5mgVyDjWmA = 32'o27745163147 ^ 32'hd40544e7;
      7'o150: EbCa5mgVyDjWmA = 32'd4139963910 ^ 32'o23524672206;
      default: EbCa5mgVyDjWmA = 32'hdead_dead;
    endcase
  end

  always_ff @(posedge clk_i) begin
    if(rst_i) begin
      parity_en <= '0;
    end
    else begin
      parity_en <= EbCa5mgVyDjWmA[32'd3951968853 ^ 32'heb8e425f];
    end
  end

  logic uJ0eNXr;

  logic [31:0] Dk3IFM518baNPDAIXFaLH;
  always_comb begin
    case ({uJ0eNXr, YAhtnxC5bxEVGCn, parity_en, Uzd, B4zEGLaAwyO6, Gdxya89mlifb})
      6'b111111: Dk3IFM518baNPDAIXFaLH = 32'o14466757122 ^ 32'h6e9ea550;
      6'd9: Dk3IFM518baNPDAIXFaLH = 32'h67e56cb ^ 32'o1416622711;
      6'h26: Dk3IFM518baNPDAIXFaLH = 32'o34711220411 ^ 32'b11101101011000000101001000001011;
      6'o25: Dk3IFM518baNPDAIXFaLH = 32'b00001111000001110101000000110111 ^ 32'b00000101010000100010001100110101;
      6'h3e: Dk3IFM518baNPDAIXFaLH = 32'h5aaabbfa ^ 32'h767d2668 ^ 32'o4644567220;
      6'd60: Dk3IFM518baNPDAIXFaLH = 32'd3272594398 ^ 32'h9bfe2a31 ^ 32'h52b48aed;
      6'h3: Dk3IFM518baNPDAIXFaLH = 32'h98e2de0d ^ 32'h92a7ad0f;
      6'o14: Dk3IFM518baNPDAIXFaLH = 32'he6591b22 ^ 32'o10543222145 ^ 32'd2844871749;
      6'h3b: Dk3IFM518baNPDAIXFaLH = 32'b01110111110101000000101001111011 ^ 32'd1226132178 ^ 32'd881079211;
      6'd44: Dk3IFM518baNPDAIXFaLH = 32'o25711406247 ^ 32'o12007662147 ^ 32'd4118551490;
      6'o67: Dk3IFM518baNPDAIXFaLH = 32'd1947992322 ^ 32'b01111110010110010111101000000000;
      6'h0: Dk3IFM518baNPDAIXFaLH = 32'o21620321142 ^ 32'h8404d160;
      6'o66: Dk3IFM518baNPDAIXFaLH = 32'o35530425455 ^ 32'o26162331047 ^ 32'b01010110111011101110101000001000;
      6'h12: Dk3IFM518baNPDAIXFaLH = 32'd456624051 ^ 32'h1e95ec2d ^ 32'd266803356;
      6'o45: Dk3IFM518baNPDAIXFaLH = 32'd1390930270 ^ 32'b01011000101000101001101001011100;
      6'd15: Dk3IFM518baNPDAIXFaLH = 32'b01110001000001001100001001101010 ^ 32'b01111011010000011011000101101000;
      6'd49: Dk3IFM518baNPDAIXFaLH = 32'o6372267241 ^ 32'o7153016643;
      6'o12: Dk3IFM518baNPDAIXFaLH = 32'b11010010100011000111111011000001 ^ 32'o33062206703;
      6'd45: Dk3IFM518baNPDAIXFaLH = 32'o11333136343 ^ 32'hb3c4159e ^ 32'o36273355177;
      6'b000101: Dk3IFM518baNPDAIXFaLH = 32'h209229e6 ^ 32'o5265655344;
      6'h3a: Dk3IFM518baNPDAIXFaLH = 32'h9cd4365b ^ 32'h96914559;
      6'h11: Dk3IFM518baNPDAIXFaLH = 32'o20271434642 ^ 32'b10001000101000110100101010100000;
      6'o15: Dk3IFM518baNPDAIXFaLH = 32'b11101000000010101100010010110111 ^ 32'o12012203035 ^ 32'b10110010011001101011000110101000;
      6'd28: Dk3IFM518baNPDAIXFaLH = 32'b00100001101110001010101010100011 ^ 32'b00101011111111011101100110100001;
      6'b101000: Dk3IFM518baNPDAIXFaLH = 32'h1b7799fd ^ 32'h1132eaff;
      6'o13: Dk3IFM518baNPDAIXFaLH = 32'h543565a5 ^ 32'o33566314175 ^ 32'o20352307332;
      6'o35: Dk3IFM518baNPDAIXFaLH = 32'o31536202452 ^ 32'b01100001100001001100010101100101 ^ 32'd2797122381;
      6'b000010: Dk3IFM518baNPDAIXFaLH = 32'o30757310151 ^ 32'b11001101111110001110001101101011;
      6'o41: Dk3IFM518baNPDAIXFaLH = 32'h84b21955 ^ 32'o21675665127;
      6'h23: Dk3IFM518baNPDAIXFaLH = 32'b00110001001000000111101011001110 ^ 32'd996477388;
      6'h6: Dk3IFM518baNPDAIXFaLH = 32'd222508838 ^ 32'b01001110011011101111111100011011 ^ 32'b01001001011010001011101100111111;
      6'h1a: Dk3IFM518baNPDAIXFaLH = 32'b11101001100011111111110010010111 ^ 32'he3ca8f95;
      6'h29: Dk3IFM518baNPDAIXFaLH = 32'b10011111011100111100111110111011 ^ 32'haecd0d8d ^ 32'o7376730464;
      6'h2e: Dk3IFM518baNPDAIXFaLH = 32'd345198075 ^ 32'o37203604521 ^ 32'd3839440808;
      6'b100010: Dk3IFM518baNPDAIXFaLH = 32'd2629307275 ^ 32'hdde50853 ^ 32'd1259892954;
      6'o30: Dk3IFM518baNPDAIXFaLH = 32'hdadceeef ^ 32'o14773635324 ^ 32'hb776a739;
      6'b101010: Dk3IFM518baNPDAIXFaLH = 32'b10110011110111110000100011010111 ^ 32'b10111001100110100111101111010101;
      6'o23: Dk3IFM518baNPDAIXFaLH = 32'he5fa5d2f ^ 32'o27067145762 ^ 32'o12730762737;
      6'd47: Dk3IFM518baNPDAIXFaLH = 32'd740697537 ^ 32'b00100110011000110101011011000011;
      6'b000100: Dk3IFM518baNPDAIXFaLH = 32'o26607741266 ^ 32'hbb73bd1b ^ 32'o712206257;
      6'o70: Dk3IFM518baNPDAIXFaLH = 32'o30653654272 ^ 32'o30276162077 ^ 32'o1604547607;
      6'he: Dk3IFM518baNPDAIXFaLH = 32'b10110000000000101111001101111001 ^ 32'b11100000111010011001100000110100 ^ 32'h5aae184f;
      6'o37: Dk3IFM518baNPDAIXFaLH = 32'o4150565566 ^ 32'b00101011111001111001000001110100;
      6'h10: Dk3IFM518baNPDAIXFaLH = 32'h810c31f0 ^ 32'h21727614 ^ 32'haa3b34e6;
      6'b110100: Dk3IFM518baNPDAIXFaLH = 32'b11011101101001001000100010111001 ^ 32'd3236754870 ^ 32'h170d0e0d;
      6'o71: Dk3IFM518baNPDAIXFaLH = 32'o26475216444 ^ 32'o17762030322 ^ 32'b11000001011110000101111011110100;
      6'o27: Dk3IFM518baNPDAIXFaLH = 32'b11000110010000000110100101101100 ^ 32'b11111110010111110101100010110000 ^ 32'b00110010010110100100101011011110;
      6'o1: Dk3IFM518baNPDAIXFaLH = 32'd4197336220 ^ 32'o1026357263 ^ 32'd4164086061;
      6'h32: Dk3IFM518baNPDAIXFaLH = 32'b00000000100110000100111010111100 ^ 32'o1267236676;
      6'h20: Dk3IFM518baNPDAIXFaLH = 32'hec49480a ^ 32'b11100110000011000011101100001000;
      6'h19: Dk3IFM518baNPDAIXFaLH = 32'h4aa9cdfb ^ 32'd3372756869 ^ 32'h89e4917c;
      6'd36: Dk3IFM518baNPDAIXFaLH = 32'b10111001011111011100010001010001 ^ 32'b10010111101100100100000010011011 ^ 32'd613087176;
      6'd48: Dk3IFM518baNPDAIXFaLH = 32'd3233831403 ^ 32'd3397724905;
      6'b110101: Dk3IFM518baNPDAIXFaLH = 32'b00110010010110100001010101001101 ^ 32'b00111000000111110110011001001111;
      6'd8: Dk3IFM518baNPDAIXFaLH = 32'b11110000011110100100000111110110 ^ 32'b11111010001111110011001011110100;
      6'd7: Dk3IFM518baNPDAIXFaLH = 32'b10001000111111011011101100000101 ^ 32'b10000010101110001100100000000111;
      6'b111101: Dk3IFM518baNPDAIXFaLH = 32'o4235655755 ^ 32'hbe95bd9a ^ 32'o22651712565;
      6'd20: Dk3IFM518baNPDAIXFaLH = 32'd1279049401 ^ 32'b01000110011110011100110110111011;
      6'b011110: Dk3IFM518baNPDAIXFaLH = 32'o6746255405 ^ 32'h56cdf100 ^ 32'd1796331783;
      6'd27: Dk3IFM518baNPDAIXFaLH = 32'd111063629 ^ 32'o34151731410 ^ 32'b11101101011111000111001001000111;
      6'o47: Dk3IFM518baNPDAIXFaLH = 32'h7889ef82 ^ 32'h1ffe37bb ^ 32'd1832037179;
      6'h16: Dk3IFM518baNPDAIXFaLH = 32'd3243279749 ^ 32'b11001011000101011111011010000111;
      6'd43: Dk3IFM518baNPDAIXFaLH = 32'd1796014351 ^ 32'h875762f5 ^ 32'o34607610370;
      6'o63: Dk3IFM518baNPDAIXFaLH = 32'b11011010110000001011011111010100 ^ 32'b11011011100010000100111110011111 ^ 32'b00001011000011011000101101001001;
      default: Dk3IFM518baNPDAIXFaLH = 32'hdead_dead;
    endcase
  end

  always_comb begin
    case ({Gdxya89mlifb, uJ0eNXr, YAhtnxC5bxEVGCn, Uzd, B4zEGLaAwyO6, lYDnXNr})
      6'h25: j22I6zJCUqZP = 32'h3dd635dc ^ 32'b00000010010011010111111111100101 ^ 32'd1977908219;
      6'o62: j22I6zJCUqZP = 32'o13611555473 ^ 32'h16b7875d ^ 32'd49180068;
      6'b010101: j22I6zJCUqZP = 32'b01111000110110011001110111000111 ^ 32'd982359434 ^ 32'd137048495;
      6'd32: j22I6zJCUqZP = 32'o27414301274 ^ 32'b00110001101001010011000111110111 ^ 32'd3354100361;
      6'o2: j22I6zJCUqZP = 32'b10100111101100010100000111110110 ^ 32'b01000110001001101111111001010111 ^ 32'd2884144739;
      6'b010110: j22I6zJCUqZP = 32'd2603225329 ^ 32'd1769493627 ^ 32'b10111000001011010111010101101000;
      6'o35: j22I6zJCUqZP = 32'o30735236007 ^ 32'h8d0a0de5;
      6'o47: j22I6zJCUqZP = 32'd2736113196 ^ 32'b11101001011010101111011111101110;
      6'd34: j22I6zJCUqZP = 32'o27055376170 ^ 32'b10010101100110110110101001110101 ^ 32'd1733404623;
      6'o23: j22I6zJCUqZP = 32'b11011011011101110100100111100100 ^ 32'd2433251366;
      6'b011011: j22I6zJCUqZP = 32'o5320022646 ^ 32'b01100001001111110001010001100100;
      6'h3: j22I6zJCUqZP = 32'h2f424ce1 ^ 32'd954329943 ^ 32'd1574737524;
      6'd35: j22I6zJCUqZP = 32'o15475635401 ^ 32'd646449859;
      6'o71: j22I6zJCUqZP = 32'b01111110010100101000101111111111 ^ 32'd875412029;
      6'o13: j22I6zJCUqZP = 32'h6049b8c4 ^ 32'o5215504406;
      6'b110111: j22I6zJCUqZP = 32'b01110110000001111111011001110010 ^ 32'd1014548400;
      6'b010001: j22I6zJCUqZP = 32'h90ac14fa ^ 32'b10011011010011111010001110110010 ^ 32'b01000001100111001000011010001010;
      6'b011100: j22I6zJCUqZP = 32'd2461837217 ^ 32'hd8c39643;
      6'o56: j22I6zJCUqZP = 32'o26446631260 ^ 32'd178967269 ^ 32'o36423550627;
      6'b111011: j22I6zJCUqZP = 32'd2875766250 ^ 32'b10001010100100110110000001100001 ^ 32'b01101011100001001110010001001001;
      6'o64: j22I6zJCUqZP = 32'o11211775022 ^ 32'd5819344;
      6'h0: j22I6zJCUqZP = 32'o6634751162 ^ 32'b00001000100111110110111100011011 ^ 32'h74938cab;
      6'd54: j22I6zJCUqZP = 32'b11101000001011000101000001110010 ^ 32'o13540451673 ^ 32'hffd1320b;
      6'o77: j22I6zJCUqZP = 32'h927b2063 ^ 32'd3851244689 ^ 32'd1032406320;
      6'd8: j22I6zJCUqZP = 32'd3635482780 ^ 32'd445641012 ^ 32'o21020350152;
      6'b001111: j22I6zJCUqZP = 32'o22226132535 ^ 32'd3626468543;
      6'o61: j22I6zJCUqZP = 32'b00111011010111001101110000100001 ^ 32'o12661302675 ^ 32'h27e6685e;
      6'd23: j22I6zJCUqZP = 32'b11010101110111010110111001010011 ^ 32'o2274551407 ^ 32'd2370866358;
      6'b000111: j22I6zJCUqZP = 32'b01100000000001101000010000111100 ^ 32'o5236332736;
      6'b000100: j22I6zJCUqZP = 32'b10011011101101000000011101111011 ^ 32'h603aded2 ^ 32'd2985420875;
      6'b101001: j22I6zJCUqZP = 32'd2123729657 ^ 32'b01001000111001001100100000010100 ^ 32'b01111100000011100111001100101111;
      6'h12: j22I6zJCUqZP = 32'b10101010000001010101101000010110 ^ 32'o13500571111 ^ 32'd3178797469;
      6'd60: j22I6zJCUqZP = 32'o1440010524 ^ 32'o14245567112 ^ 32'h2469cedc;
      6'd56: j22I6zJCUqZP = 32'hf3ae5e17 ^ 32'b10110001100110111100001111101010 ^ 32'b00001000010010101010110000111111;
      6'd5: j22I6zJCUqZP = 32'd2683208167 ^ 32'o32544330005;
      6'b010100: j22I6zJCUqZP = 32'b11100001001000111110001111010011 ^ 32'h9677cafc ^ 32'o7512614315;
      6'b011111: j22I6zJCUqZP = 32'hea2aadf9 ^ 32'b10100000010101011001110000011011;
      6'h19: j22I6zJCUqZP = 32'o23534443314 ^ 32'hd70d770e;
      6'd45: j22I6zJCUqZP = 32'd979130504 ^ 32'o27762533332 ^ 32'o31772357620;
      6'b101010: j22I6zJCUqZP = 32'b11100100011101000101001100011101 ^ 32'o25602661337;
      6'b001110: j22I6zJCUqZP = 32'h56167a48 ^ 32'b01001001001000001101100110111010 ^ 32'h55499210;
      6'o1: j22I6zJCUqZP = 32'b11110101101001000001000111110011 ^ 32'b10111111110110110010000000110001;
      6'b101100: j22I6zJCUqZP = 32'd284674992 ^ 32'b01010110010010110110000000010000 ^ 32'o1460715142;
      6'h6: j22I6zJCUqZP = 32'o765222175 ^ 32'd1302992287;
      6'h28: j22I6zJCUqZP = 32'hd944ecc1 ^ 32'h4501e378 ^ 32'b11010110001110100011111001111011;
      6'h10: j22I6zJCUqZP = 32'h9cb44fb1 ^ 32'b10110000011001011010001001011101 ^ 32'b01100110101011101101110000101110;
      6'd13: j22I6zJCUqZP = 32'd3601912019 ^ 32'o23463760461;
      6'o12: j22I6zJCUqZP = 32'b11101111111111111101101011111110 ^ 32'ha580eb3c;
      6'o65: j22I6zJCUqZP = 32'hcb0e052f ^ 32'd729170173 ^ 32'o25201672020;
      6'h3e: j22I6zJCUqZP = 32'hb95893f5 ^ 32'o14442637462 ^ 32'd2544672005;
      6'd47: j22I6zJCUqZP = 32'd2219559306 ^ 32'd3459577928;
      6'o44: j22I6zJCUqZP = 32'd1789602431 ^ 32'b00100000110101000001101110111101;
      6'b100110: j22I6zJCUqZP = 32'hfacb78bd ^ 32'heb2d6c32 ^ 32'h5b99254d;
      6'b111010: j22I6zJCUqZP = 32'b10101100010110110100010101111111 ^ 32'b11100110001001000111010010111101;
      6'd48: j22I6zJCUqZP = 32'd1913282486 ^ 32'o7035267164;
      6'o30: j22I6zJCUqZP = 32'b11100101011101000001010100001001 ^ 32'b10101111000010110010010011001011;
      6'd51: j22I6zJCUqZP = 32'o12312441473 ^ 32'h182d5a25 ^ 32'o136024334;
      6'b011010: j22I6zJCUqZP = 32'o13074315357 ^ 32'h128eab2d;
      6'b001001: j22I6zJCUqZP = 32'b11101110011111111111111011011010 ^ 32'o24400147430;
      6'b011110: j22I6zJCUqZP = 32'b11111010000101100000001000010010 ^ 32'd1096486261 ^ 32'hf1323e85;
      6'd61: j22I6zJCUqZP = 32'b00110111110010010011101001101001 ^ 32'd2109082539;
      6'b001100: j22I6zJCUqZP = 32'd3808382059 ^ 32'hfecff04f ^ 32'h564f8dc6;
      6'd43: j22I6zJCUqZP = 32'b10100100000000001000001000100001 ^ 32'd4001346531;
      6'd33: j22I6zJCUqZP = 32'o24751310673 ^ 32'o1374711003 ^ 32'he629327a;
      default: j22I6zJCUqZP = 32'hdead_dead;
    endcase
  end

  assign uJ0eNXr = (Y2pd == (32'd1189161525 ^ 32'o1460235663 ^ 32'o11210010622));
  logic [31:0] uNUkwrQnCG;
  always_comb begin
    case ({YAhtnxC5bxEVGCn, parity_en, busy, Gdxya89mlifb, uJ0eNXr, Uzd})
      6'b011101: uNUkwrQnCG = 32'o26720515475 ^ 32'he16cbe92 ^ 32'o11061734725;
      6'b000010: uNUkwrQnCG = 32'd3437905050 ^ 32'd1777622794 ^ 32'hbbf787ea;
      6'b110111: uNUkwrQnCG = 32'd3633841046 ^ 32'haa601fcd ^ 32'd1813086497;
      6'o1: uNUkwrQnCG = 32'o3362340612 ^ 32'b00000101001000000101110111110000;
      6'o51: uNUkwrQnCG = 32'b10101011110111011000011100010101 ^ 32'hb5341b6f;
      6'h1c: uNUkwrQnCG = 32'o15007305301 ^ 32'b10100110011000011100001001100010 ^ 32'hd095d4d9;
      6'b101011: uNUkwrQnCG = 32'o17402511660 ^ 32'b01100100011010000011011000010110 ^ 32'b00000110100010110011100111011100;
      6'o37: uNUkwrQnCG = 32'b10101101111110011100111011011011 ^ 32'o26304051641;
      6'o14: uNUkwrQnCG = 32'b00011001000101111011111110001100 ^ 32'b00000111111111100010001111110110;
      6'b111100: uNUkwrQnCG = 32'd592909713 ^ 32'd1035897323;
      6'b100011: uNUkwrQnCG = 32'b00011111100000101110100101001111 ^ 32'd23819573;
      6'h17: uNUkwrQnCG = 32'd3849944139 ^ 32'd4220576049;
      6'd4: uNUkwrQnCG = 32'o34360106777 ^ 32'hfd291185;
      6'b110010: uNUkwrQnCG = 32'd1294144214 ^ 32'd4083829118 ^ 32'b10100000101000001100011111010010;
      6'b100000: uNUkwrQnCG = 32'hd94ed3ca ^ 32'h9c1237e5 ^ 32'h5bb57855;
      6'd34: uNUkwrQnCG = 32'o35613471603 ^ 32'h77edf0e ^ 32'o36756230367;
      6'h34: uNUkwrQnCG = 32'h2dae2ae ^ 32'b11011110111011011001000101000000 ^ 32'o30267567624;
      6'b110000: uNUkwrQnCG = 32'b01101101001110110001001110010111 ^ 32'o16364507755;
      6'o24: uNUkwrQnCG = 32'd269181137 ^ 32'o3241056357 ^ 32'h1466a044;
      6'd16: uNUkwrQnCG = 32'd1581802107 ^ 32'd1084358145;
      6'o46: uNUkwrQnCG = 32'h2368c922 ^ 32'd3127744844 ^ 32'b10000111111011001100110000010100;
      6'o36: uNUkwrQnCG = 32'd3630626997 ^ 32'd396194741 ^ 32'd3507623802;
      6'd15: uNUkwrQnCG = 32'ha7e7ad7b ^ 32'hb90e3001;
      6'b001101: uNUkwrQnCG = 32'b11101101000000011000000100010100 ^ 32'b11110011111010000001110101101110;
      6'o75: uNUkwrQnCG = 32'hf76eb2c3 ^ 32'o7076534461 ^ 32'd3514668936;
      6'd11: uNUkwrQnCG = 32'b10010010100100000011001100010000 ^ 32'ha13521fe ^ 32'o5523107224;
      6'd27: uNUkwrQnCG = 32'he895aa8b ^ 32'b01001011101001011001110000011110 ^ 32'b10111101110110011010101011101111;
      6'b010011: uNUkwrQnCG = 32'd2624686312 ^ 32'o20246012222;
      6'd63: uNUkwrQnCG = 32'o26532705111 ^ 32'b01111100100000001011101101101001 ^ 32'hd702ac5a;
      6'd57: uNUkwrQnCG = 32'o2356375073 ^ 32'o4417675522 ^ 32'h296f1d13;
      6'b011000: uNUkwrQnCG = 32'b00001001011110110110101101000111 ^ 32'b00010111100100101111011100111101;
      6'h3e: uNUkwrQnCG = 32'b00010010010110011010010001011110 ^ 32'h28f2c8d6 ^ 32'd608366834;
      6'o72: uNUkwrQnCG = 32'd794064492 ^ 32'd1118138119 ^ 32'd1930986769;
      6'd46: uNUkwrQnCG = 32'd1131470182 ^ 32'b11011110111101100110001101011001 ^ 32'b10000011011011110010001001000101;
      6'o26: uNUkwrQnCG = 32'b10101001110001011000110100110100 ^ 32'hb72c114e;
      6'd36: uNUkwrQnCG = 32'h33a6199e ^ 32'd3736286497 ^ 32'hf3fcb0c5;
      6'd6: uNUkwrQnCG = 32'd983123423 ^ 32'o4434154645;
      6'b000111: uNUkwrQnCG = 32'hd304af81 ^ 32'o34330761122 ^ 32'b00101110100011101101000010101001;
      6'b101010: uNUkwrQnCG = 32'd1263231941 ^ 32'd1436745663;
      6'o12: uNUkwrQnCG = 32'h5f4f3849 ^ 32'b01000001101001101010010000110011;
      6'h3b: uNUkwrQnCG = 32'b11001010010011110011110110011101 ^ 32'hd4a6a1e7;
      6'h0: uNUkwrQnCG = 32'b11000101110111111001010011101010 ^ 32'd3677751440;
      6'h2f: uNUkwrQnCG = 32'd3757892785 ^ 32'd3239410123;
      6'b110011: uNUkwrQnCG = 32'h841fb21 ^ 32'o22222142124 ^ 32'h84e0a30f;
      6'o22: uNUkwrQnCG = 32'h907e649d ^ 32'h8e97f8e7;
      6'd37: uNUkwrQnCG = 32'b10110011011010001000101000110000 ^ 32'o25540213112;
      6'h11: uNUkwrQnCG = 32'o23750123616 ^ 32'd3620524801 ^ 32'o12641364365;
      6'b101100: uNUkwrQnCG = 32'b10010100110000000111001010101010 ^ 32'b10001010001010011110111011010000;
      6'o11: uNUkwrQnCG = 32'h7e7044b4 ^ 32'b01100000100110011101100011001110;
      6'b110110: uNUkwrQnCG = 32'd1841593561 ^ 32'o16313360243;
      6'd25: uNUkwrQnCG = 32'o12212375610 ^ 32'b01001100110000000110011111110010;
      6'o50: uNUkwrQnCG = 32'b01111110110111110101000010011101 ^ 32'b01100000001101101100110011100111;
      6'b101101: uNUkwrQnCG = 32'o7131252100 ^ 32'h278cc83a;
      6'h3: uNUkwrQnCG = 32'b10011000100010110011000101101010 ^ 32'o20630526420;
      6'd5: uNUkwrQnCG = 32'hb3a10773 ^ 32'd3420061772 ^ 32'b01100110100100101001101101000101;
      6'o65: uNUkwrQnCG = 32'b11001110110011101000100000100010 ^ 32'o5343050031 ^ 32'b11111011101010110100010001000001;
      6'd56: uNUkwrQnCG = 32'h1f151683 ^ 32'h1fc8af9;
      6'o47: uNUkwrQnCG = 32'hb08bfd31 ^ 32'b00111001101111110011101111010010 ^ 32'h97dd5b99;
      6'h31: uNUkwrQnCG = 32'd1348320380 ^ 32'b11110010101010011101110001111110 ^ 32'hbc1dfc78;
      6'd26: uNUkwrQnCG = 32'o5234755557 ^ 32'h349a4715;
      6'h8: uNUkwrQnCG = 32'o35527417352 ^ 32'd304754521 ^ 32'he19dadc9;
      6'd33: uNUkwrQnCG = 32'o772510167 ^ 32'h6c9c8ee2 ^ 32'h759f82ef;
      6'h15: uNUkwrQnCG = 32'd2503373721 ^ 32'h27f9407c ^ 32'o25411527637;
      6'd14: uNUkwrQnCG = 32'hc76d7c0d ^ 32'b11011001100001001110000001110111;
      default: uNUkwrQnCG = 32'hdead_dead;
    endcase
  end
  logic [1:0] Ab1IpiFqqV2O;
  assign Ab1IpiFqqV2O = ra2VgcBEzc[1:0];

  always_ff @(posedge clk_i) begin
    if(rst_i) begin
      stopbit <= 1;
    end
    else if (Dk3IFM518baNPDAIXFaLH[32'h6cc8350c ^ 32'hfebafa7c ^ 32'h9272cf7b]) begin
      stopbit <= 2'b01;
    end
    else if(uNUkwrQnCG[32'hdf990339 ^ 32'o6234265624 ^ 32'o35572064245]) begin
      stopbit <= Ab1IpiFqqV2O;
    end
    else begin
      stopbit <= stopbit;
    end
  end

  logic [31:0] CQSw5rojmDCtLn8X9U8DKok;

  always_ff @(posedge clk_i) begin
    if(rst_i) begin
      eCNnNC8kn <= 32'hc5fb985e ^ 32'o20537213333 ^ 32'h40868e85;
    end
    else if (CQSw5rojmDCtLn8X9U8DKok[32'o33214101136 ^ 32'hda308244]) begin
      eCNnNC8kn <= 32'ha7944dfa ^ 32'd983050913 ^ 32'b10011101000011000110011101011011;
    end
    else if(j22I6zJCUqZP[32'b11010110110101111110111010110001 ^ 32'd3604475572]) begin
      case(Y2pd)
        32'd2718025493 ^ 32'hcd5ebaa6 ^ 32'd1868529075: eCNnNC8kn <= data;
        32'b10110000000000100111100101110010 ^ 32'b10000110010010011110001101100010 ^ 32'o6622715034: eCNnNC8kn <= baudrate;
        32'hf60c972b ^ 32'b11110010000011011011001110100010 ^ 32'b00000100000000010010010010000001: eCNnNC8kn <= busy;
        32'hec292561 ^ 32'h82ef4211 ^ 32'd1858496356: eCNnNC8kn <= stopbit;
        32'd1889123409 ^ 32'b00011010100100111001111000101111 ^ 32'b01101010000010100010001001101110: eCNnNC8kn <= parity_en;
        default: eCNnNC8kn <= eCNnNC8kn;
      endcase
    end
    else begin
      eCNnNC8kn <= eCNnNC8kn;
    end
  end
  always_comb begin
    case ({Gdxya89mlifb, uJ0eNXr, YAhtnxC5bxEVGCn, Uzd, B4zEGLaAwyO6, lYDnXNr})
      6'h5: CQSw5rojmDCtLn8X9U8DKok = 32'd2033132964 ^ 32'o2340302472;
      6'd26: CQSw5rojmDCtLn8X9U8DKok = 32'h11ea89c9 ^ 32'd2068064599;
      6'h2: CQSw5rojmDCtLn8X9U8DKok = 32'he7522c70 ^ 32'd3238617996 ^ 32'd1291186018;
      6'b100001: CQSw5rojmDCtLn8X9U8DKok = 32'd197517268 ^ 32'b01100001011010110111111101001010;
      6'h33: CQSw5rojmDCtLn8X9U8DKok = 32'b01011100000000101001001111111011 ^ 32'd917255013;
      6'h29: CQSw5rojmDCtLn8X9U8DKok = 32'd2025856909 ^ 32'b00000011100100000101011010000110 ^ 32'o2177564625;
      6'h13: CQSw5rojmDCtLn8X9U8DKok = 32'o754213012 ^ 32'd1830794900;
      6'o34: CQSw5rojmDCtLn8X9U8DKok = 32'b01110010101000001000111111010101 ^ 32'b00011000000011100010111101001011;
      6'd35: CQSw5rojmDCtLn8X9U8DKok = 32'b10110001000101000000010001111000 ^ 32'hdbbaa4e6;
      6'o10: CQSw5rojmDCtLn8X9U8DKok = 32'd2603620176 ^ 32'd4272611475 ^ 32'o1715053535;
      6'b001101: CQSw5rojmDCtLn8X9U8DKok = 32'b11101001110010011001100111110011 ^ 32'h8367396d;
      6'h14: CQSw5rojmDCtLn8X9U8DKok = 32'o21372505664 ^ 32'hd4d3f128 ^ 32'd899144194;
      6'o50: CQSw5rojmDCtLn8X9U8DKok = 32'b01110001110101101001100011100100 ^ 32'b00011011011110000011100001111010;
      6'b001011: CQSw5rojmDCtLn8X9U8DKok = 32'hd6af009c ^ 32'hbc01a002;
      6'b101111: CQSw5rojmDCtLn8X9U8DKok = 32'b10010011001000101000000001100101 ^ 32'b11111101100011000010000011111011;
      6'b011000: CQSw5rojmDCtLn8X9U8DKok = 32'd501010915 ^ 32'd2003988861;
      6'h30: CQSw5rojmDCtLn8X9U8DKok = 32'b01101000010101010010111111110001 ^ 32'o4617237654 ^ 32'd617001155;
      6'b000110: CQSw5rojmDCtLn8X9U8DKok = 32'h8a528e00 ^ 32'b01110001110111010101101000101000 ^ 32'b10010001001000010111010010110110;
      6'b100000: CQSw5rojmDCtLn8X9U8DKok = 32'o10362123012 ^ 32'd364343967 ^ 32'h3cd1740b;
      6'b100110: CQSw5rojmDCtLn8X9U8DKok = 32'hb154cbc4 ^ 32'b11011011111110100110101101011010;
      6'o53: CQSw5rojmDCtLn8X9U8DKok = 32'b11100101001010011010011100001111 ^ 32'd3469954698 ^ 32'd1096042779;
      6'd10: CQSw5rojmDCtLn8X9U8DKok = 32'd244763119 ^ 32'o35533106523 ^ 32'b10001001010101001110010000100010;
      6'h3: CQSw5rojmDCtLn8X9U8DKok = 32'o2701541250 ^ 32'h7da86236;
      6'b111001: CQSw5rojmDCtLn8X9U8DKok = 32'b01111000011011010001100111100100 ^ 32'o2260734572;
      6'b010101: CQSw5rojmDCtLn8X9U8DKok = 32'b10111000010100001011010111001011 ^ 32'd3822284759 ^ 32'o6113275202;
      6'd61: CQSw5rojmDCtLn8X9U8DKok = 32'd337875502 ^ 32'o26013577235 ^ 32'b11001110101000111100110000101101;
      6'd12: CQSw5rojmDCtLn8X9U8DKok = 32'b01000011111010111000010101100111 ^ 32'hc204e65f ^ 32'd3946955686;
      6'h32: CQSw5rojmDCtLn8X9U8DKok = 32'hda520725 ^ 32'b10110000111111001010011110111011;
      6'b100101: CQSw5rojmDCtLn8X9U8DKok = 32'd2503901057 ^ 32'hff90df1f;
      6'h27: CQSw5rojmDCtLn8X9U8DKok = 32'b00010011110100111010001110001111 ^ 32'h797d0311;
      6'd23: CQSw5rojmDCtLn8X9U8DKok = 32'd1075940450 ^ 32'd3592570192 ^ 32'b11111100101011010110100110101100;
      6'o4: CQSw5rojmDCtLn8X9U8DKok = 32'hb8939f3c ^ 32'hd23d3fa2;
      6'h34: CQSw5rojmDCtLn8X9U8DKok = 32'b01111001011011100000111001001010 ^ 32'h13c0aed4;
      6'd27: CQSw5rojmDCtLn8X9U8DKok = 32'b11010100000101110010001000100100 ^ 32'b10111110101110011000001010111010;
      6'hf: CQSw5rojmDCtLn8X9U8DKok = 32'b01110111110111001001000001000000 ^ 32'd494022878;
      6'o7: CQSw5rojmDCtLn8X9U8DKok = 32'd1615240095 ^ 32'o27534222440 ^ 32'b10110111100110010001111000100001;
      6'o73: CQSw5rojmDCtLn8X9U8DKok = 32'd755412675 ^ 32'b00101100101000001110111110010000 ^ 32'b01101011000010001110000111001101;
      6'b111111: CQSw5rojmDCtLn8X9U8DKok = 32'b11011000001110101010010111001111 ^ 32'hb6940551;
      6'h35: CQSw5rojmDCtLn8X9U8DKok = 32'd547625192 ^ 32'h4a0ab876;
      6'b010010: CQSw5rojmDCtLn8X9U8DKok = 32'd683123692 ^ 32'o10206201562;
      6'b011110: CQSw5rojmDCtLn8X9U8DKok = 32'o10147360137 ^ 32'o23002312075 ^ 32'b10110011001110101101010011111100;
      6'o0: CQSw5rojmDCtLn8X9U8DKok = 32'h5481f694 ^ 32'o7613653012;
      6'h9: CQSw5rojmDCtLn8X9U8DKok = 32'd2144664520 ^ 32'b10011011110011010000110010010011 ^ 32'd2394380229;
      6'd29: CQSw5rojmDCtLn8X9U8DKok = 32'b10010001000110101000111111011001 ^ 32'o37355027507;
      6'o31: CQSw5rojmDCtLn8X9U8DKok = 32'o23674052347 ^ 32'hf45ef479;
      6'd45: CQSw5rojmDCtLn8X9U8DKok = 32'b11111111000110001101100110001111 ^ 32'h6591f6de ^ 32'b11110000001001111000111111001111;
      6'o56: CQSw5rojmDCtLn8X9U8DKok = 32'o37732425536 ^ 32'o13045422624 ^ 32'hc952ae54;
      6'b110111: CQSw5rojmDCtLn8X9U8DKok = 32'o37776403363 ^ 32'd2505352813;
      6'h10: CQSw5rojmDCtLn8X9U8DKok = 32'o13525330336 ^ 32'h4922df44 ^ 32'd2128203524;
      6'b010001: CQSw5rojmDCtLn8X9U8DKok = 32'd3122673693 ^ 32'h4c079be7 ^ 32'b10011100100010010000001101100100;
      6'o61: CQSw5rojmDCtLn8X9U8DKok = 32'h1fc89785 ^ 32'b01110101011001100011011100011011;
      6'b010110: CQSw5rojmDCtLn8X9U8DKok = 32'd1628030088 ^ 32'hba76416;
      6'b101010: CQSw5rojmDCtLn8X9U8DKok = 32'h6a9ddddf ^ 32'h337d41;
      6'h1: CQSw5rojmDCtLn8X9U8DKok = 32'd1387559939 ^ 32'b01000011010110001010101110010111 ^ 32'h7b42770a;
      6'd58: CQSw5rojmDCtLn8X9U8DKok = 32'd2089823772 ^ 32'h3048a8e2 ^ 32'h26762660;
      6'b111100: CQSw5rojmDCtLn8X9U8DKok = 32'o4756252415 ^ 32'o12612402221 ^ 32'o3317370402;
      6'd14: CQSw5rojmDCtLn8X9U8DKok = 32'd182870714 ^ 32'o14022141044;
      6'h24: CQSw5rojmDCtLn8X9U8DKok = 32'o25666657060 ^ 32'o2666633564 ^ 32'o32253544732;
      6'd56: CQSw5rojmDCtLn8X9U8DKok = 32'h75de70f6 ^ 32'd527487080;
      6'd31: CQSw5rojmDCtLn8X9U8DKok = 32'o6113143612 ^ 32'o25574455561 ^ 32'hf6703c65;
      6'd34: CQSw5rojmDCtLn8X9U8DKok = 32'o23751047343 ^ 32'o15307350572 ^ 32'h9e173f07;
      6'd62: CQSw5rojmDCtLn8X9U8DKok = 32'b11000000100110110011100011010101 ^ 32'd31920334 ^ 32'hafd28885;
      6'd44: CQSw5rojmDCtLn8X9U8DKok = 32'd1378007252 ^ 32'd948705354;
      6'b110110: CQSw5rojmDCtLn8X9U8DKok = 32'b01101100100010001111010100011001 ^ 32'd45723561 ^ 32'h49ffa2e;
      default: CQSw5rojmDCtLn8X9U8DKok = 32'hdead_dead;
    endcase
  end

  assign tzBmaC = (Y2pd == (32'b01010111001110010000000010100100 ^ 32'o10727355447 ^ 32'h1064db8f));
endmodule
